module IOB(
  input  [31:0] io_in_0,
  output [31:0] io_out_0
);
  assign io_out_0 = io_in_0; // @[IOB.scala 53:42]
endmodule
module Muxn(
  input         io_config,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  output [31:0] io_out
);
  assign io_out = io_config ? io_in_1 : io_in_0; // @[Multiplexer.scala 20:10]
endmodule
module ConfigMem(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [31:0] io_cfg_data,
  output        io_out_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg  regs_0; // @[ConfigMem.scala 27:21]
  assign io_out_0 = regs_0; // @[ConfigMem.scala 52:45]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  regs_0 = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      regs_0 <= 1'h0;
    end else if (io_cfg_en) begin
      regs_0 <= io_cfg_data[0];
    end
  end
endmodule
module IOB_16(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  output [31:0] io_out_0
);
  wire  Muxn_io_config; // @[IOB.scala 36:41]
  wire [31:0] Muxn_io_in_0; // @[IOB.scala 36:41]
  wire [31:0] Muxn_io_in_1; // @[IOB.scala 36:41]
  wire [31:0] Muxn_io_out; // @[IOB.scala 36:41]
  wire  ConfigMem_clock; // @[IOB.scala 37:21]
  wire  ConfigMem_reset; // @[IOB.scala 37:21]
  wire  ConfigMem_io_cfg_en; // @[IOB.scala 37:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[IOB.scala 37:21]
  wire  ConfigMem_io_out_0; // @[IOB.scala 37:21]
  wire  _T_1 = 10'ha == io_cfg_addr[11:2]; // @[IOB.scala 38:50]
  Muxn Muxn ( // @[IOB.scala 36:41]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_out(Muxn_io_out)
  );
  ConfigMem ConfigMem ( // @[IOB.scala 37:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  assign io_out_0 = Muxn_io_out; // @[IOB.scala 48:17]
  assign Muxn_io_config = ConfigMem_io_out_0; // @[IOB.scala 49:22]
  assign Muxn_io_in_0 = io_in_0; // @[IOB.scala 46:23]
  assign Muxn_io_in_1 = io_in_1; // @[IOB.scala 46:23]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[IOB.scala 38:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[IOB.scala 40:21]
endmodule
module IOB_17(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  output [31:0] io_out_0
);
  wire  Muxn_io_config; // @[IOB.scala 36:41]
  wire [31:0] Muxn_io_in_0; // @[IOB.scala 36:41]
  wire [31:0] Muxn_io_in_1; // @[IOB.scala 36:41]
  wire [31:0] Muxn_io_out; // @[IOB.scala 36:41]
  wire  ConfigMem_clock; // @[IOB.scala 37:21]
  wire  ConfigMem_reset; // @[IOB.scala 37:21]
  wire  ConfigMem_io_cfg_en; // @[IOB.scala 37:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[IOB.scala 37:21]
  wire  ConfigMem_io_out_0; // @[IOB.scala 37:21]
  wire  _T_1 = 10'hb == io_cfg_addr[11:2]; // @[IOB.scala 38:50]
  Muxn Muxn ( // @[IOB.scala 36:41]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_out(Muxn_io_out)
  );
  ConfigMem ConfigMem ( // @[IOB.scala 37:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  assign io_out_0 = Muxn_io_out; // @[IOB.scala 48:17]
  assign Muxn_io_config = ConfigMem_io_out_0; // @[IOB.scala 49:22]
  assign Muxn_io_in_0 = io_in_0; // @[IOB.scala 46:23]
  assign Muxn_io_in_1 = io_in_1; // @[IOB.scala 46:23]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[IOB.scala 38:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[IOB.scala 40:21]
endmodule
module IOB_18(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  output [31:0] io_out_0
);
  wire  Muxn_io_config; // @[IOB.scala 36:41]
  wire [31:0] Muxn_io_in_0; // @[IOB.scala 36:41]
  wire [31:0] Muxn_io_in_1; // @[IOB.scala 36:41]
  wire [31:0] Muxn_io_out; // @[IOB.scala 36:41]
  wire  ConfigMem_clock; // @[IOB.scala 37:21]
  wire  ConfigMem_reset; // @[IOB.scala 37:21]
  wire  ConfigMem_io_cfg_en; // @[IOB.scala 37:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[IOB.scala 37:21]
  wire  ConfigMem_io_out_0; // @[IOB.scala 37:21]
  wire  _T_1 = 10'hc == io_cfg_addr[11:2]; // @[IOB.scala 38:50]
  Muxn Muxn ( // @[IOB.scala 36:41]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_out(Muxn_io_out)
  );
  ConfigMem ConfigMem ( // @[IOB.scala 37:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  assign io_out_0 = Muxn_io_out; // @[IOB.scala 48:17]
  assign Muxn_io_config = ConfigMem_io_out_0; // @[IOB.scala 49:22]
  assign Muxn_io_in_0 = io_in_0; // @[IOB.scala 46:23]
  assign Muxn_io_in_1 = io_in_1; // @[IOB.scala 46:23]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[IOB.scala 38:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[IOB.scala 40:21]
endmodule
module IOB_19(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  output [31:0] io_out_0
);
  wire  Muxn_io_config; // @[IOB.scala 36:41]
  wire [31:0] Muxn_io_in_0; // @[IOB.scala 36:41]
  wire [31:0] Muxn_io_in_1; // @[IOB.scala 36:41]
  wire [31:0] Muxn_io_out; // @[IOB.scala 36:41]
  wire  ConfigMem_clock; // @[IOB.scala 37:21]
  wire  ConfigMem_reset; // @[IOB.scala 37:21]
  wire  ConfigMem_io_cfg_en; // @[IOB.scala 37:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[IOB.scala 37:21]
  wire  ConfigMem_io_out_0; // @[IOB.scala 37:21]
  wire  _T_1 = 10'hd == io_cfg_addr[11:2]; // @[IOB.scala 38:50]
  Muxn Muxn ( // @[IOB.scala 36:41]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_out(Muxn_io_out)
  );
  ConfigMem ConfigMem ( // @[IOB.scala 37:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  assign io_out_0 = Muxn_io_out; // @[IOB.scala 48:17]
  assign Muxn_io_config = ConfigMem_io_out_0; // @[IOB.scala 49:22]
  assign Muxn_io_in_0 = io_in_0; // @[IOB.scala 46:23]
  assign Muxn_io_in_1 = io_in_1; // @[IOB.scala 46:23]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[IOB.scala 38:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[IOB.scala 40:21]
endmodule
module IOB_20(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  output [31:0] io_out_0
);
  wire  Muxn_io_config; // @[IOB.scala 36:41]
  wire [31:0] Muxn_io_in_0; // @[IOB.scala 36:41]
  wire [31:0] Muxn_io_in_1; // @[IOB.scala 36:41]
  wire [31:0] Muxn_io_out; // @[IOB.scala 36:41]
  wire  ConfigMem_clock; // @[IOB.scala 37:21]
  wire  ConfigMem_reset; // @[IOB.scala 37:21]
  wire  ConfigMem_io_cfg_en; // @[IOB.scala 37:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[IOB.scala 37:21]
  wire  ConfigMem_io_out_0; // @[IOB.scala 37:21]
  wire  _T_1 = 10'he == io_cfg_addr[11:2]; // @[IOB.scala 38:50]
  Muxn Muxn ( // @[IOB.scala 36:41]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_out(Muxn_io_out)
  );
  ConfigMem ConfigMem ( // @[IOB.scala 37:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  assign io_out_0 = Muxn_io_out; // @[IOB.scala 48:17]
  assign Muxn_io_config = ConfigMem_io_out_0; // @[IOB.scala 49:22]
  assign Muxn_io_in_0 = io_in_0; // @[IOB.scala 46:23]
  assign Muxn_io_in_1 = io_in_1; // @[IOB.scala 46:23]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[IOB.scala 38:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[IOB.scala 40:21]
endmodule
module IOB_21(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  output [31:0] io_out_0
);
  wire  Muxn_io_config; // @[IOB.scala 36:41]
  wire [31:0] Muxn_io_in_0; // @[IOB.scala 36:41]
  wire [31:0] Muxn_io_in_1; // @[IOB.scala 36:41]
  wire [31:0] Muxn_io_out; // @[IOB.scala 36:41]
  wire  ConfigMem_clock; // @[IOB.scala 37:21]
  wire  ConfigMem_reset; // @[IOB.scala 37:21]
  wire  ConfigMem_io_cfg_en; // @[IOB.scala 37:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[IOB.scala 37:21]
  wire  ConfigMem_io_out_0; // @[IOB.scala 37:21]
  wire  _T_1 = 10'hf == io_cfg_addr[11:2]; // @[IOB.scala 38:50]
  Muxn Muxn ( // @[IOB.scala 36:41]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_out(Muxn_io_out)
  );
  ConfigMem ConfigMem ( // @[IOB.scala 37:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  assign io_out_0 = Muxn_io_out; // @[IOB.scala 48:17]
  assign Muxn_io_config = ConfigMem_io_out_0; // @[IOB.scala 49:22]
  assign Muxn_io_in_0 = io_in_0; // @[IOB.scala 46:23]
  assign Muxn_io_in_1 = io_in_1; // @[IOB.scala 46:23]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[IOB.scala 38:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[IOB.scala 40:21]
endmodule
module IOB_22(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  output [31:0] io_out_0
);
  wire  Muxn_io_config; // @[IOB.scala 36:41]
  wire [31:0] Muxn_io_in_0; // @[IOB.scala 36:41]
  wire [31:0] Muxn_io_in_1; // @[IOB.scala 36:41]
  wire [31:0] Muxn_io_out; // @[IOB.scala 36:41]
  wire  ConfigMem_clock; // @[IOB.scala 37:21]
  wire  ConfigMem_reset; // @[IOB.scala 37:21]
  wire  ConfigMem_io_cfg_en; // @[IOB.scala 37:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[IOB.scala 37:21]
  wire  ConfigMem_io_out_0; // @[IOB.scala 37:21]
  wire  _T_1 = 10'h10 == io_cfg_addr[11:2]; // @[IOB.scala 38:50]
  Muxn Muxn ( // @[IOB.scala 36:41]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_out(Muxn_io_out)
  );
  ConfigMem ConfigMem ( // @[IOB.scala 37:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  assign io_out_0 = Muxn_io_out; // @[IOB.scala 48:17]
  assign Muxn_io_config = ConfigMem_io_out_0; // @[IOB.scala 49:22]
  assign Muxn_io_in_0 = io_in_0; // @[IOB.scala 46:23]
  assign Muxn_io_in_1 = io_in_1; // @[IOB.scala 46:23]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[IOB.scala 38:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[IOB.scala 40:21]
endmodule
module IOB_23(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  output [31:0] io_out_0
);
  wire  Muxn_io_config; // @[IOB.scala 36:41]
  wire [31:0] Muxn_io_in_0; // @[IOB.scala 36:41]
  wire [31:0] Muxn_io_in_1; // @[IOB.scala 36:41]
  wire [31:0] Muxn_io_out; // @[IOB.scala 36:41]
  wire  ConfigMem_clock; // @[IOB.scala 37:21]
  wire  ConfigMem_reset; // @[IOB.scala 37:21]
  wire  ConfigMem_io_cfg_en; // @[IOB.scala 37:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[IOB.scala 37:21]
  wire  ConfigMem_io_out_0; // @[IOB.scala 37:21]
  wire  _T_1 = 10'h11 == io_cfg_addr[11:2]; // @[IOB.scala 38:50]
  Muxn Muxn ( // @[IOB.scala 36:41]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_out(Muxn_io_out)
  );
  ConfigMem ConfigMem ( // @[IOB.scala 37:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  assign io_out_0 = Muxn_io_out; // @[IOB.scala 48:17]
  assign Muxn_io_config = ConfigMem_io_out_0; // @[IOB.scala 49:22]
  assign Muxn_io_in_0 = io_in_0; // @[IOB.scala 46:23]
  assign Muxn_io_in_1 = io_in_1; // @[IOB.scala 46:23]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[IOB.scala 38:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[IOB.scala 40:21]
endmodule
module IOB_24(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  output [31:0] io_out_0
);
  wire  Muxn_io_config; // @[IOB.scala 36:41]
  wire [31:0] Muxn_io_in_0; // @[IOB.scala 36:41]
  wire [31:0] Muxn_io_in_1; // @[IOB.scala 36:41]
  wire [31:0] Muxn_io_out; // @[IOB.scala 36:41]
  wire  ConfigMem_clock; // @[IOB.scala 37:21]
  wire  ConfigMem_reset; // @[IOB.scala 37:21]
  wire  ConfigMem_io_cfg_en; // @[IOB.scala 37:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[IOB.scala 37:21]
  wire  ConfigMem_io_out_0; // @[IOB.scala 37:21]
  wire  _T_1 = 10'hb5 == io_cfg_addr[11:2]; // @[IOB.scala 38:50]
  Muxn Muxn ( // @[IOB.scala 36:41]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_out(Muxn_io_out)
  );
  ConfigMem ConfigMem ( // @[IOB.scala 37:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  assign io_out_0 = Muxn_io_out; // @[IOB.scala 48:17]
  assign Muxn_io_config = ConfigMem_io_out_0; // @[IOB.scala 49:22]
  assign Muxn_io_in_0 = io_in_0; // @[IOB.scala 46:23]
  assign Muxn_io_in_1 = io_in_1; // @[IOB.scala 46:23]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[IOB.scala 38:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[IOB.scala 40:21]
endmodule
module IOB_25(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  output [31:0] io_out_0
);
  wire  Muxn_io_config; // @[IOB.scala 36:41]
  wire [31:0] Muxn_io_in_0; // @[IOB.scala 36:41]
  wire [31:0] Muxn_io_in_1; // @[IOB.scala 36:41]
  wire [31:0] Muxn_io_out; // @[IOB.scala 36:41]
  wire  ConfigMem_clock; // @[IOB.scala 37:21]
  wire  ConfigMem_reset; // @[IOB.scala 37:21]
  wire  ConfigMem_io_cfg_en; // @[IOB.scala 37:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[IOB.scala 37:21]
  wire  ConfigMem_io_out_0; // @[IOB.scala 37:21]
  wire  _T_1 = 10'hb6 == io_cfg_addr[11:2]; // @[IOB.scala 38:50]
  Muxn Muxn ( // @[IOB.scala 36:41]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_out(Muxn_io_out)
  );
  ConfigMem ConfigMem ( // @[IOB.scala 37:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  assign io_out_0 = Muxn_io_out; // @[IOB.scala 48:17]
  assign Muxn_io_config = ConfigMem_io_out_0; // @[IOB.scala 49:22]
  assign Muxn_io_in_0 = io_in_0; // @[IOB.scala 46:23]
  assign Muxn_io_in_1 = io_in_1; // @[IOB.scala 46:23]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[IOB.scala 38:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[IOB.scala 40:21]
endmodule
module IOB_26(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  output [31:0] io_out_0
);
  wire  Muxn_io_config; // @[IOB.scala 36:41]
  wire [31:0] Muxn_io_in_0; // @[IOB.scala 36:41]
  wire [31:0] Muxn_io_in_1; // @[IOB.scala 36:41]
  wire [31:0] Muxn_io_out; // @[IOB.scala 36:41]
  wire  ConfigMem_clock; // @[IOB.scala 37:21]
  wire  ConfigMem_reset; // @[IOB.scala 37:21]
  wire  ConfigMem_io_cfg_en; // @[IOB.scala 37:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[IOB.scala 37:21]
  wire  ConfigMem_io_out_0; // @[IOB.scala 37:21]
  wire  _T_1 = 10'hb7 == io_cfg_addr[11:2]; // @[IOB.scala 38:50]
  Muxn Muxn ( // @[IOB.scala 36:41]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_out(Muxn_io_out)
  );
  ConfigMem ConfigMem ( // @[IOB.scala 37:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  assign io_out_0 = Muxn_io_out; // @[IOB.scala 48:17]
  assign Muxn_io_config = ConfigMem_io_out_0; // @[IOB.scala 49:22]
  assign Muxn_io_in_0 = io_in_0; // @[IOB.scala 46:23]
  assign Muxn_io_in_1 = io_in_1; // @[IOB.scala 46:23]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[IOB.scala 38:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[IOB.scala 40:21]
endmodule
module IOB_27(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  output [31:0] io_out_0
);
  wire  Muxn_io_config; // @[IOB.scala 36:41]
  wire [31:0] Muxn_io_in_0; // @[IOB.scala 36:41]
  wire [31:0] Muxn_io_in_1; // @[IOB.scala 36:41]
  wire [31:0] Muxn_io_out; // @[IOB.scala 36:41]
  wire  ConfigMem_clock; // @[IOB.scala 37:21]
  wire  ConfigMem_reset; // @[IOB.scala 37:21]
  wire  ConfigMem_io_cfg_en; // @[IOB.scala 37:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[IOB.scala 37:21]
  wire  ConfigMem_io_out_0; // @[IOB.scala 37:21]
  wire  _T_1 = 10'hb8 == io_cfg_addr[11:2]; // @[IOB.scala 38:50]
  Muxn Muxn ( // @[IOB.scala 36:41]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_out(Muxn_io_out)
  );
  ConfigMem ConfigMem ( // @[IOB.scala 37:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  assign io_out_0 = Muxn_io_out; // @[IOB.scala 48:17]
  assign Muxn_io_config = ConfigMem_io_out_0; // @[IOB.scala 49:22]
  assign Muxn_io_in_0 = io_in_0; // @[IOB.scala 46:23]
  assign Muxn_io_in_1 = io_in_1; // @[IOB.scala 46:23]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[IOB.scala 38:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[IOB.scala 40:21]
endmodule
module IOB_28(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  output [31:0] io_out_0
);
  wire  Muxn_io_config; // @[IOB.scala 36:41]
  wire [31:0] Muxn_io_in_0; // @[IOB.scala 36:41]
  wire [31:0] Muxn_io_in_1; // @[IOB.scala 36:41]
  wire [31:0] Muxn_io_out; // @[IOB.scala 36:41]
  wire  ConfigMem_clock; // @[IOB.scala 37:21]
  wire  ConfigMem_reset; // @[IOB.scala 37:21]
  wire  ConfigMem_io_cfg_en; // @[IOB.scala 37:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[IOB.scala 37:21]
  wire  ConfigMem_io_out_0; // @[IOB.scala 37:21]
  wire  _T_1 = 10'hb9 == io_cfg_addr[11:2]; // @[IOB.scala 38:50]
  Muxn Muxn ( // @[IOB.scala 36:41]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_out(Muxn_io_out)
  );
  ConfigMem ConfigMem ( // @[IOB.scala 37:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  assign io_out_0 = Muxn_io_out; // @[IOB.scala 48:17]
  assign Muxn_io_config = ConfigMem_io_out_0; // @[IOB.scala 49:22]
  assign Muxn_io_in_0 = io_in_0; // @[IOB.scala 46:23]
  assign Muxn_io_in_1 = io_in_1; // @[IOB.scala 46:23]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[IOB.scala 38:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[IOB.scala 40:21]
endmodule
module IOB_29(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  output [31:0] io_out_0
);
  wire  Muxn_io_config; // @[IOB.scala 36:41]
  wire [31:0] Muxn_io_in_0; // @[IOB.scala 36:41]
  wire [31:0] Muxn_io_in_1; // @[IOB.scala 36:41]
  wire [31:0] Muxn_io_out; // @[IOB.scala 36:41]
  wire  ConfigMem_clock; // @[IOB.scala 37:21]
  wire  ConfigMem_reset; // @[IOB.scala 37:21]
  wire  ConfigMem_io_cfg_en; // @[IOB.scala 37:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[IOB.scala 37:21]
  wire  ConfigMem_io_out_0; // @[IOB.scala 37:21]
  wire  _T_1 = 10'hba == io_cfg_addr[11:2]; // @[IOB.scala 38:50]
  Muxn Muxn ( // @[IOB.scala 36:41]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_out(Muxn_io_out)
  );
  ConfigMem ConfigMem ( // @[IOB.scala 37:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  assign io_out_0 = Muxn_io_out; // @[IOB.scala 48:17]
  assign Muxn_io_config = ConfigMem_io_out_0; // @[IOB.scala 49:22]
  assign Muxn_io_in_0 = io_in_0; // @[IOB.scala 46:23]
  assign Muxn_io_in_1 = io_in_1; // @[IOB.scala 46:23]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[IOB.scala 38:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[IOB.scala 40:21]
endmodule
module IOB_30(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  output [31:0] io_out_0
);
  wire  Muxn_io_config; // @[IOB.scala 36:41]
  wire [31:0] Muxn_io_in_0; // @[IOB.scala 36:41]
  wire [31:0] Muxn_io_in_1; // @[IOB.scala 36:41]
  wire [31:0] Muxn_io_out; // @[IOB.scala 36:41]
  wire  ConfigMem_clock; // @[IOB.scala 37:21]
  wire  ConfigMem_reset; // @[IOB.scala 37:21]
  wire  ConfigMem_io_cfg_en; // @[IOB.scala 37:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[IOB.scala 37:21]
  wire  ConfigMem_io_out_0; // @[IOB.scala 37:21]
  wire  _T_1 = 10'hbb == io_cfg_addr[11:2]; // @[IOB.scala 38:50]
  Muxn Muxn ( // @[IOB.scala 36:41]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_out(Muxn_io_out)
  );
  ConfigMem ConfigMem ( // @[IOB.scala 37:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  assign io_out_0 = Muxn_io_out; // @[IOB.scala 48:17]
  assign Muxn_io_config = ConfigMem_io_out_0; // @[IOB.scala 49:22]
  assign Muxn_io_in_0 = io_in_0; // @[IOB.scala 46:23]
  assign Muxn_io_in_1 = io_in_1; // @[IOB.scala 46:23]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[IOB.scala 38:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[IOB.scala 40:21]
endmodule
module IOB_31(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  output [31:0] io_out_0
);
  wire  Muxn_io_config; // @[IOB.scala 36:41]
  wire [31:0] Muxn_io_in_0; // @[IOB.scala 36:41]
  wire [31:0] Muxn_io_in_1; // @[IOB.scala 36:41]
  wire [31:0] Muxn_io_out; // @[IOB.scala 36:41]
  wire  ConfigMem_clock; // @[IOB.scala 37:21]
  wire  ConfigMem_reset; // @[IOB.scala 37:21]
  wire  ConfigMem_io_cfg_en; // @[IOB.scala 37:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[IOB.scala 37:21]
  wire  ConfigMem_io_out_0; // @[IOB.scala 37:21]
  wire  _T_1 = 10'hbc == io_cfg_addr[11:2]; // @[IOB.scala 38:50]
  Muxn Muxn ( // @[IOB.scala 36:41]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_out(Muxn_io_out)
  );
  ConfigMem ConfigMem ( // @[IOB.scala 37:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  assign io_out_0 = Muxn_io_out; // @[IOB.scala 48:17]
  assign Muxn_io_config = ConfigMem_io_out_0; // @[IOB.scala 49:22]
  assign Muxn_io_in_0 = io_in_0; // @[IOB.scala 46:23]
  assign Muxn_io_in_1 = io_in_1; // @[IOB.scala 46:23]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[IOB.scala 38:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[IOB.scala 40:21]
endmodule
module ALU(
  input  [3:0]  io_config,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  output [31:0] io_out
);
  wire [31:0] _T_4 = io_in_0 + io_in_1; // @[Operations.scala 124:41]
  wire [31:0] _T_8 = io_in_0 - io_in_1; // @[Operations.scala 126:41]
  wire [63:0] _T_11 = io_in_0 * io_in_1; // @[Operations.scala 128:41]
  wire [31:0] _T_14 = io_in_0 & io_in_1; // @[Operations.scala 138:41]
  wire [31:0] _T_17 = io_in_0 | io_in_1; // @[Operations.scala 140:41]
  wire [31:0] _T_20 = io_in_0 ^ io_in_1; // @[Operations.scala 142:41]
  wire  _T_21 = 4'h0 == io_config; // @[Mux.scala 80:60]
  wire [31:0] _T_22 = _T_21 ? io_in_0 : 32'h0; // @[Mux.scala 80:57]
  wire  _T_23 = 4'h1 == io_config; // @[Mux.scala 80:60]
  wire [31:0] _T_24 = _T_23 ? _T_4 : _T_22; // @[Mux.scala 80:57]
  wire  _T_25 = 4'h2 == io_config; // @[Mux.scala 80:60]
  wire [31:0] _T_26 = _T_25 ? _T_8 : _T_24; // @[Mux.scala 80:57]
  wire  _T_27 = 4'h3 == io_config; // @[Mux.scala 80:60]
  wire [63:0] _T_28 = _T_27 ? _T_11 : {{32'd0}, _T_26}; // @[Mux.scala 80:57]
  wire  _T_29 = 4'h4 == io_config; // @[Mux.scala 80:60]
  wire [63:0] _T_30 = _T_29 ? {{32'd0}, _T_14} : _T_28; // @[Mux.scala 80:57]
  wire  _T_31 = 4'h5 == io_config; // @[Mux.scala 80:60]
  wire [63:0] _T_32 = _T_31 ? {{32'd0}, _T_17} : _T_30; // @[Mux.scala 80:57]
  wire  _T_33 = 4'h6 == io_config; // @[Mux.scala 80:60]
  wire [63:0] _T_34 = _T_33 ? {{32'd0}, _T_20} : _T_32; // @[Mux.scala 80:57]
  assign io_out = _T_34[31:0]; // @[ALU.scala 25:10]
endmodule
module RF(
  input         clock,
  input         reset,
  input         io_en,
  input  [31:0] io_in_0,
  output [31:0] io_out_0,
  output [31:0] io_out_1
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] regs_0; // @[RegFile.scala 24:21]
  assign io_out_0 = regs_0; // @[RegFile.scala 37:42]
  assign io_out_1 = regs_0; // @[RegFile.scala 37:42]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  regs_0 = _RAND_0[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      regs_0 <= 32'h0;
    end else if (io_en) begin
      regs_0 <= io_in_0;
    end
  end
endmodule
module DelayPipe(
  input         clock,
  input         reset,
  input         io_en,
  input  [2:0]  io_config,
  input  [31:0] io_in,
  output [31:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] regs_0; // @[DelayPipe.scala 22:21]
  reg [31:0] regs_1; // @[DelayPipe.scala 22:21]
  reg [31:0] regs_2; // @[DelayPipe.scala 22:21]
  reg [31:0] regs_3; // @[DelayPipe.scala 22:21]
  reg [31:0] regs_4; // @[DelayPipe.scala 22:21]
  reg [2:0] wptr; // @[DelayPipe.scala 23:21]
  reg [2:0] rptr; // @[DelayPipe.scala 24:21]
  wire  _T_1 = wptr < 3'h4; // @[DelayPipe.scala 26:23]
  wire  _T_2 = io_en & _T_1; // @[DelayPipe.scala 26:14]
  wire [2:0] _T_4 = wptr + 3'h1; // @[DelayPipe.scala 27:17]
  wire  _T_7 = _T_4 >= io_config; // @[DelayPipe.scala 32:17]
  wire [2:0] _T_11 = _T_4 - io_config; // @[DelayPipe.scala 33:24]
  wire [2:0] _T_13 = 3'h6 + wptr; // @[DelayPipe.scala 35:30]
  wire [2:0] _T_15 = _T_13 - io_config; // @[DelayPipe.scala 35:37]
  wire  _T_16 = io_config > 3'h0; // @[DelayPipe.scala 39:28]
  wire  _T_17 = io_en & _T_16; // @[DelayPipe.scala 39:14]
  reg [2:0] cnt; // @[DelayPipe.scala 43:20]
  wire  _T_18 = ~io_en; // @[DelayPipe.scala 44:8]
  wire  _T_19 = cnt < io_config; // @[DelayPipe.scala 46:18]
  wire [2:0] _T_21 = cnt + 3'h1; // @[DelayPipe.scala 47:16]
  wire  _T_22 = 3'h0 == io_config; // @[DelayPipe.scala 50:22]
  wire  _T_23 = io_en & _T_22; // @[DelayPipe.scala 50:14]
  wire  _T_24 = cnt == io_config; // @[DelayPipe.scala 52:28]
  wire  _T_25 = io_en & _T_24; // @[DelayPipe.scala 52:20]
  wire [31:0] _GEN_15 = 3'h1 == rptr ? regs_1 : regs_0; // @[DelayPipe.scala 53:12]
  wire [31:0] _GEN_16 = 3'h2 == rptr ? regs_2 : _GEN_15; // @[DelayPipe.scala 53:12]
  wire [31:0] _GEN_17 = 3'h3 == rptr ? regs_3 : _GEN_16; // @[DelayPipe.scala 53:12]
  wire [31:0] _GEN_18 = 3'h4 == rptr ? regs_4 : _GEN_17; // @[DelayPipe.scala 53:12]
  wire [31:0] _GEN_19 = _T_25 ? _GEN_18 : 32'h0; // @[DelayPipe.scala 52:43]
  assign io_out = _T_23 ? io_in : _GEN_19; // @[DelayPipe.scala 51:12 DelayPipe.scala 53:12 DelayPipe.scala 55:12]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  regs_0 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  regs_1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  regs_2 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  regs_3 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  regs_4 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  wptr = _RAND_5[2:0];
  _RAND_6 = {1{`RANDOM}};
  rptr = _RAND_6[2:0];
  _RAND_7 = {1{`RANDOM}};
  cnt = _RAND_7[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      regs_0 <= 32'h0;
    end else if (_T_17) begin
      if (3'h0 == wptr) begin
        regs_0 <= io_in;
      end
    end
    if (reset) begin
      regs_1 <= 32'h0;
    end else if (_T_17) begin
      if (3'h1 == wptr) begin
        regs_1 <= io_in;
      end
    end
    if (reset) begin
      regs_2 <= 32'h0;
    end else if (_T_17) begin
      if (3'h2 == wptr) begin
        regs_2 <= io_in;
      end
    end
    if (reset) begin
      regs_3 <= 32'h0;
    end else if (_T_17) begin
      if (3'h3 == wptr) begin
        regs_3 <= io_in;
      end
    end
    if (reset) begin
      regs_4 <= 32'h0;
    end else if (_T_17) begin
      if (3'h4 == wptr) begin
        regs_4 <= io_in;
      end
    end
    if (reset) begin
      wptr <= 3'h0;
    end else if (_T_2) begin
      wptr <= _T_4;
    end else begin
      wptr <= 3'h0;
    end
    if (reset) begin
      rptr <= 3'h0;
    end else if (_T_7) begin
      rptr <= _T_11;
    end else begin
      rptr <= _T_15;
    end
    if (reset) begin
      cnt <= 3'h0;
    end else if (_T_18) begin
      cnt <= 3'h0;
    end else if (_T_19) begin
      cnt <= _T_21;
    end
  end
endmodule
module Muxn_16(
  input  [2:0]  io_config,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  output [31:0] io_out
);
  wire  _T_2 = 3'h1 == io_config; // @[Mux.scala 80:60]
  wire [31:0] _T_3 = _T_2 ? io_in_1 : io_in_0; // @[Mux.scala 80:57]
  wire  _T_4 = 3'h2 == io_config; // @[Mux.scala 80:60]
  wire [31:0] _T_5 = _T_4 ? io_in_2 : _T_3; // @[Mux.scala 80:57]
  wire  _T_6 = 3'h3 == io_config; // @[Mux.scala 80:60]
  wire [31:0] _T_7 = _T_6 ? io_in_3 : _T_5; // @[Mux.scala 80:57]
  wire  _T_8 = 3'h4 == io_config; // @[Mux.scala 80:60]
  wire [31:0] _T_9 = _T_8 ? io_in_4 : _T_7; // @[Mux.scala 80:57]
  wire  _T_10 = 3'h5 == io_config; // @[Mux.scala 80:60]
  assign io_out = _T_10 ? io_in_5 : _T_9; // @[Multiplexer.scala 20:10]
endmodule
module ConfigMem_16(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input         io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [47:0] io_out_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [47:0] regs_0; // @[ConfigMem.scala 27:21]
  wire  _T_1 = ~io_cfg_addr; // @[ConfigMem.scala 39:38]
  wire  _T_2 = io_cfg_en & _T_1; // @[ConfigMem.scala 39:22]
  wire [47:0] _T_4 = {regs_0[47:32],io_cfg_data}; // @[Cat.scala 29:58]
  wire [47:0] _GEN_0 = _T_2 ? _T_4 : regs_0; // @[ConfigMem.scala 39:47]
  wire  _T_6 = io_cfg_en & io_cfg_addr; // @[ConfigMem.scala 39:22]
  wire [63:0] _T_8 = {io_cfg_data,regs_0[31:0]}; // @[Cat.scala 29:58]
  wire [63:0] _GEN_1 = _T_6 ? _T_8 : {{16'd0}, _GEN_0}; // @[ConfigMem.scala 39:47]
  assign io_out_0 = regs_0; // @[ConfigMem.scala 52:45]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  regs_0 = _RAND_0[47:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      regs_0 <= 48'h0;
    end else begin
      regs_0 <= _GEN_1[47:0];
    end
  end
endmodule
module GPE(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [3:0] alu_io_config; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 50:19]
  wire [31:0] alu_io_out; // @[PE.scala 50:19]
  wire  rf_clock; // @[PE.scala 51:18]
  wire  rf_reset; // @[PE.scala 51:18]
  wire  rf_io_en; // @[PE.scala 51:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 51:18]
  wire  DelayPipe_clock; // @[PE.scala 52:54]
  wire  DelayPipe_reset; // @[PE.scala 52:54]
  wire  DelayPipe_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 52:54]
  wire  DelayPipe_1_clock; // @[PE.scala 52:54]
  wire  DelayPipe_1_reset; // @[PE.scala 52:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 52:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 55:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 55:49]
  wire  cfg_clock; // @[PE.scala 89:19]
  wire  cfg_reset; // @[PE.scala 89:19]
  wire  cfg_io_cfg_en; // @[PE.scala 89:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 89:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 89:19]
  wire [47:0] cfg_io_out_0; // @[PE.scala 89:19]
  wire  _T_1 = 10'h1c == io_cfg_addr[11:2]; // @[PE.scala 90:48]
  wire [47:0] cfgOut = cfg_io_out_0; // @[PE.scala 96:20 PE.scala 97:10]
  ALU alu ( // @[PE.scala 50:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 51:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 52:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 52:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_16 Muxn ( // @[PE.scala 55:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_16 Muxn_1 ( // @[PE.scala 55:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_16 cfg ( // @[PE.scala 89:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 77:13]
  assign alu_io_config = cfgOut[35:32]; // @[PE.scala 100:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 71:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 71:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 75:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 76:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_io_config = cfgOut[38:36]; // @[PE.scala 113:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 70:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_1_io_config = cfgOut[41:39]; // @[PE.scala 113:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 70:23]
  assign Muxn_io_config = cfgOut[44:42]; // @[PE.scala 121:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 62:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 62:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 62:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 62:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign Muxn_1_io_config = cfgOut[47:45]; // @[PE.scala 121:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 62:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 62:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 62:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 62:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 90:17]
  assign cfg_io_cfg_addr = io_cfg_addr[0]; // @[PE.scala 91:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 92:19]
endmodule
module GPE_1(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [3:0] alu_io_config; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 50:19]
  wire [31:0] alu_io_out; // @[PE.scala 50:19]
  wire  rf_clock; // @[PE.scala 51:18]
  wire  rf_reset; // @[PE.scala 51:18]
  wire  rf_io_en; // @[PE.scala 51:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 51:18]
  wire  DelayPipe_clock; // @[PE.scala 52:54]
  wire  DelayPipe_reset; // @[PE.scala 52:54]
  wire  DelayPipe_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 52:54]
  wire  DelayPipe_1_clock; // @[PE.scala 52:54]
  wire  DelayPipe_1_reset; // @[PE.scala 52:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 52:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 55:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 55:49]
  wire  cfg_clock; // @[PE.scala 89:19]
  wire  cfg_reset; // @[PE.scala 89:19]
  wire  cfg_io_cfg_en; // @[PE.scala 89:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 89:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 89:19]
  wire [47:0] cfg_io_out_0; // @[PE.scala 89:19]
  wire  _T_1 = 10'h1d == io_cfg_addr[11:2]; // @[PE.scala 90:48]
  wire [47:0] cfgOut = cfg_io_out_0; // @[PE.scala 96:20 PE.scala 97:10]
  ALU alu ( // @[PE.scala 50:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 51:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 52:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 52:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_16 Muxn ( // @[PE.scala 55:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_16 Muxn_1 ( // @[PE.scala 55:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_16 cfg ( // @[PE.scala 89:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 77:13]
  assign alu_io_config = cfgOut[35:32]; // @[PE.scala 100:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 71:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 71:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 75:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 76:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_io_config = cfgOut[38:36]; // @[PE.scala 113:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 70:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_1_io_config = cfgOut[41:39]; // @[PE.scala 113:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 70:23]
  assign Muxn_io_config = cfgOut[44:42]; // @[PE.scala 121:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 62:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 62:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 62:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 62:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign Muxn_1_io_config = cfgOut[47:45]; // @[PE.scala 121:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 62:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 62:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 62:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 62:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 90:17]
  assign cfg_io_cfg_addr = io_cfg_addr[0]; // @[PE.scala 91:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 92:19]
endmodule
module GPE_2(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [3:0] alu_io_config; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 50:19]
  wire [31:0] alu_io_out; // @[PE.scala 50:19]
  wire  rf_clock; // @[PE.scala 51:18]
  wire  rf_reset; // @[PE.scala 51:18]
  wire  rf_io_en; // @[PE.scala 51:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 51:18]
  wire  DelayPipe_clock; // @[PE.scala 52:54]
  wire  DelayPipe_reset; // @[PE.scala 52:54]
  wire  DelayPipe_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 52:54]
  wire  DelayPipe_1_clock; // @[PE.scala 52:54]
  wire  DelayPipe_1_reset; // @[PE.scala 52:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 52:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 55:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 55:49]
  wire  cfg_clock; // @[PE.scala 89:19]
  wire  cfg_reset; // @[PE.scala 89:19]
  wire  cfg_io_cfg_en; // @[PE.scala 89:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 89:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 89:19]
  wire [47:0] cfg_io_out_0; // @[PE.scala 89:19]
  wire  _T_1 = 10'h1e == io_cfg_addr[11:2]; // @[PE.scala 90:48]
  wire [47:0] cfgOut = cfg_io_out_0; // @[PE.scala 96:20 PE.scala 97:10]
  ALU alu ( // @[PE.scala 50:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 51:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 52:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 52:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_16 Muxn ( // @[PE.scala 55:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_16 Muxn_1 ( // @[PE.scala 55:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_16 cfg ( // @[PE.scala 89:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 77:13]
  assign alu_io_config = cfgOut[35:32]; // @[PE.scala 100:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 71:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 71:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 75:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 76:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_io_config = cfgOut[38:36]; // @[PE.scala 113:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 70:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_1_io_config = cfgOut[41:39]; // @[PE.scala 113:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 70:23]
  assign Muxn_io_config = cfgOut[44:42]; // @[PE.scala 121:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 62:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 62:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 62:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 62:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign Muxn_1_io_config = cfgOut[47:45]; // @[PE.scala 121:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 62:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 62:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 62:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 62:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 90:17]
  assign cfg_io_cfg_addr = io_cfg_addr[0]; // @[PE.scala 91:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 92:19]
endmodule
module GPE_3(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [3:0] alu_io_config; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 50:19]
  wire [31:0] alu_io_out; // @[PE.scala 50:19]
  wire  rf_clock; // @[PE.scala 51:18]
  wire  rf_reset; // @[PE.scala 51:18]
  wire  rf_io_en; // @[PE.scala 51:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 51:18]
  wire  DelayPipe_clock; // @[PE.scala 52:54]
  wire  DelayPipe_reset; // @[PE.scala 52:54]
  wire  DelayPipe_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 52:54]
  wire  DelayPipe_1_clock; // @[PE.scala 52:54]
  wire  DelayPipe_1_reset; // @[PE.scala 52:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 52:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 55:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 55:49]
  wire  cfg_clock; // @[PE.scala 89:19]
  wire  cfg_reset; // @[PE.scala 89:19]
  wire  cfg_io_cfg_en; // @[PE.scala 89:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 89:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 89:19]
  wire [47:0] cfg_io_out_0; // @[PE.scala 89:19]
  wire  _T_1 = 10'h1f == io_cfg_addr[11:2]; // @[PE.scala 90:48]
  wire [47:0] cfgOut = cfg_io_out_0; // @[PE.scala 96:20 PE.scala 97:10]
  ALU alu ( // @[PE.scala 50:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 51:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 52:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 52:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_16 Muxn ( // @[PE.scala 55:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_16 Muxn_1 ( // @[PE.scala 55:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_16 cfg ( // @[PE.scala 89:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 77:13]
  assign alu_io_config = cfgOut[35:32]; // @[PE.scala 100:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 71:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 71:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 75:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 76:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_io_config = cfgOut[38:36]; // @[PE.scala 113:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 70:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_1_io_config = cfgOut[41:39]; // @[PE.scala 113:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 70:23]
  assign Muxn_io_config = cfgOut[44:42]; // @[PE.scala 121:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 62:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 62:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 62:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 62:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign Muxn_1_io_config = cfgOut[47:45]; // @[PE.scala 121:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 62:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 62:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 62:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 62:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 90:17]
  assign cfg_io_cfg_addr = io_cfg_addr[0]; // @[PE.scala 91:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 92:19]
endmodule
module GPE_4(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [3:0] alu_io_config; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 50:19]
  wire [31:0] alu_io_out; // @[PE.scala 50:19]
  wire  rf_clock; // @[PE.scala 51:18]
  wire  rf_reset; // @[PE.scala 51:18]
  wire  rf_io_en; // @[PE.scala 51:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 51:18]
  wire  DelayPipe_clock; // @[PE.scala 52:54]
  wire  DelayPipe_reset; // @[PE.scala 52:54]
  wire  DelayPipe_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 52:54]
  wire  DelayPipe_1_clock; // @[PE.scala 52:54]
  wire  DelayPipe_1_reset; // @[PE.scala 52:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 52:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 55:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 55:49]
  wire  cfg_clock; // @[PE.scala 89:19]
  wire  cfg_reset; // @[PE.scala 89:19]
  wire  cfg_io_cfg_en; // @[PE.scala 89:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 89:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 89:19]
  wire [47:0] cfg_io_out_0; // @[PE.scala 89:19]
  wire  _T_1 = 10'h20 == io_cfg_addr[11:2]; // @[PE.scala 90:48]
  wire [47:0] cfgOut = cfg_io_out_0; // @[PE.scala 96:20 PE.scala 97:10]
  ALU alu ( // @[PE.scala 50:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 51:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 52:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 52:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_16 Muxn ( // @[PE.scala 55:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_16 Muxn_1 ( // @[PE.scala 55:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_16 cfg ( // @[PE.scala 89:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 77:13]
  assign alu_io_config = cfgOut[35:32]; // @[PE.scala 100:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 71:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 71:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 75:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 76:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_io_config = cfgOut[38:36]; // @[PE.scala 113:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 70:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_1_io_config = cfgOut[41:39]; // @[PE.scala 113:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 70:23]
  assign Muxn_io_config = cfgOut[44:42]; // @[PE.scala 121:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 62:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 62:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 62:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 62:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign Muxn_1_io_config = cfgOut[47:45]; // @[PE.scala 121:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 62:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 62:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 62:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 62:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 90:17]
  assign cfg_io_cfg_addr = io_cfg_addr[0]; // @[PE.scala 91:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 92:19]
endmodule
module GPE_5(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [3:0] alu_io_config; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 50:19]
  wire [31:0] alu_io_out; // @[PE.scala 50:19]
  wire  rf_clock; // @[PE.scala 51:18]
  wire  rf_reset; // @[PE.scala 51:18]
  wire  rf_io_en; // @[PE.scala 51:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 51:18]
  wire  DelayPipe_clock; // @[PE.scala 52:54]
  wire  DelayPipe_reset; // @[PE.scala 52:54]
  wire  DelayPipe_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 52:54]
  wire  DelayPipe_1_clock; // @[PE.scala 52:54]
  wire  DelayPipe_1_reset; // @[PE.scala 52:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 52:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 55:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 55:49]
  wire  cfg_clock; // @[PE.scala 89:19]
  wire  cfg_reset; // @[PE.scala 89:19]
  wire  cfg_io_cfg_en; // @[PE.scala 89:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 89:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 89:19]
  wire [47:0] cfg_io_out_0; // @[PE.scala 89:19]
  wire  _T_1 = 10'h21 == io_cfg_addr[11:2]; // @[PE.scala 90:48]
  wire [47:0] cfgOut = cfg_io_out_0; // @[PE.scala 96:20 PE.scala 97:10]
  ALU alu ( // @[PE.scala 50:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 51:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 52:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 52:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_16 Muxn ( // @[PE.scala 55:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_16 Muxn_1 ( // @[PE.scala 55:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_16 cfg ( // @[PE.scala 89:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 77:13]
  assign alu_io_config = cfgOut[35:32]; // @[PE.scala 100:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 71:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 71:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 75:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 76:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_io_config = cfgOut[38:36]; // @[PE.scala 113:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 70:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_1_io_config = cfgOut[41:39]; // @[PE.scala 113:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 70:23]
  assign Muxn_io_config = cfgOut[44:42]; // @[PE.scala 121:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 62:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 62:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 62:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 62:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign Muxn_1_io_config = cfgOut[47:45]; // @[PE.scala 121:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 62:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 62:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 62:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 62:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 90:17]
  assign cfg_io_cfg_addr = io_cfg_addr[0]; // @[PE.scala 91:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 92:19]
endmodule
module GPE_6(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [3:0] alu_io_config; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 50:19]
  wire [31:0] alu_io_out; // @[PE.scala 50:19]
  wire  rf_clock; // @[PE.scala 51:18]
  wire  rf_reset; // @[PE.scala 51:18]
  wire  rf_io_en; // @[PE.scala 51:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 51:18]
  wire  DelayPipe_clock; // @[PE.scala 52:54]
  wire  DelayPipe_reset; // @[PE.scala 52:54]
  wire  DelayPipe_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 52:54]
  wire  DelayPipe_1_clock; // @[PE.scala 52:54]
  wire  DelayPipe_1_reset; // @[PE.scala 52:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 52:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 55:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 55:49]
  wire  cfg_clock; // @[PE.scala 89:19]
  wire  cfg_reset; // @[PE.scala 89:19]
  wire  cfg_io_cfg_en; // @[PE.scala 89:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 89:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 89:19]
  wire [47:0] cfg_io_out_0; // @[PE.scala 89:19]
  wire  _T_1 = 10'h22 == io_cfg_addr[11:2]; // @[PE.scala 90:48]
  wire [47:0] cfgOut = cfg_io_out_0; // @[PE.scala 96:20 PE.scala 97:10]
  ALU alu ( // @[PE.scala 50:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 51:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 52:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 52:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_16 Muxn ( // @[PE.scala 55:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_16 Muxn_1 ( // @[PE.scala 55:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_16 cfg ( // @[PE.scala 89:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 77:13]
  assign alu_io_config = cfgOut[35:32]; // @[PE.scala 100:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 71:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 71:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 75:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 76:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_io_config = cfgOut[38:36]; // @[PE.scala 113:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 70:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_1_io_config = cfgOut[41:39]; // @[PE.scala 113:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 70:23]
  assign Muxn_io_config = cfgOut[44:42]; // @[PE.scala 121:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 62:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 62:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 62:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 62:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign Muxn_1_io_config = cfgOut[47:45]; // @[PE.scala 121:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 62:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 62:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 62:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 62:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 90:17]
  assign cfg_io_cfg_addr = io_cfg_addr[0]; // @[PE.scala 91:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 92:19]
endmodule
module GPE_7(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [3:0] alu_io_config; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 50:19]
  wire [31:0] alu_io_out; // @[PE.scala 50:19]
  wire  rf_clock; // @[PE.scala 51:18]
  wire  rf_reset; // @[PE.scala 51:18]
  wire  rf_io_en; // @[PE.scala 51:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 51:18]
  wire  DelayPipe_clock; // @[PE.scala 52:54]
  wire  DelayPipe_reset; // @[PE.scala 52:54]
  wire  DelayPipe_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 52:54]
  wire  DelayPipe_1_clock; // @[PE.scala 52:54]
  wire  DelayPipe_1_reset; // @[PE.scala 52:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 52:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 55:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 55:49]
  wire  cfg_clock; // @[PE.scala 89:19]
  wire  cfg_reset; // @[PE.scala 89:19]
  wire  cfg_io_cfg_en; // @[PE.scala 89:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 89:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 89:19]
  wire [47:0] cfg_io_out_0; // @[PE.scala 89:19]
  wire  _T_1 = 10'h23 == io_cfg_addr[11:2]; // @[PE.scala 90:48]
  wire [47:0] cfgOut = cfg_io_out_0; // @[PE.scala 96:20 PE.scala 97:10]
  ALU alu ( // @[PE.scala 50:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 51:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 52:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 52:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_16 Muxn ( // @[PE.scala 55:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_16 Muxn_1 ( // @[PE.scala 55:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_16 cfg ( // @[PE.scala 89:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 77:13]
  assign alu_io_config = cfgOut[35:32]; // @[PE.scala 100:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 71:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 71:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 75:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 76:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_io_config = cfgOut[38:36]; // @[PE.scala 113:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 70:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_1_io_config = cfgOut[41:39]; // @[PE.scala 113:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 70:23]
  assign Muxn_io_config = cfgOut[44:42]; // @[PE.scala 121:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 62:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 62:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 62:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 62:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign Muxn_1_io_config = cfgOut[47:45]; // @[PE.scala 121:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 62:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 62:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 62:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 62:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 90:17]
  assign cfg_io_cfg_addr = io_cfg_addr[0]; // @[PE.scala 91:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 92:19]
endmodule
module GPE_8(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [3:0] alu_io_config; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 50:19]
  wire [31:0] alu_io_out; // @[PE.scala 50:19]
  wire  rf_clock; // @[PE.scala 51:18]
  wire  rf_reset; // @[PE.scala 51:18]
  wire  rf_io_en; // @[PE.scala 51:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 51:18]
  wire  DelayPipe_clock; // @[PE.scala 52:54]
  wire  DelayPipe_reset; // @[PE.scala 52:54]
  wire  DelayPipe_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 52:54]
  wire  DelayPipe_1_clock; // @[PE.scala 52:54]
  wire  DelayPipe_1_reset; // @[PE.scala 52:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 52:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 55:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 55:49]
  wire  cfg_clock; // @[PE.scala 89:19]
  wire  cfg_reset; // @[PE.scala 89:19]
  wire  cfg_io_cfg_en; // @[PE.scala 89:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 89:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 89:19]
  wire [47:0] cfg_io_out_0; // @[PE.scala 89:19]
  wire  _T_1 = 10'h2e == io_cfg_addr[11:2]; // @[PE.scala 90:48]
  wire [47:0] cfgOut = cfg_io_out_0; // @[PE.scala 96:20 PE.scala 97:10]
  ALU alu ( // @[PE.scala 50:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 51:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 52:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 52:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_16 Muxn ( // @[PE.scala 55:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_16 Muxn_1 ( // @[PE.scala 55:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_16 cfg ( // @[PE.scala 89:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 77:13]
  assign alu_io_config = cfgOut[35:32]; // @[PE.scala 100:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 71:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 71:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 75:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 76:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_io_config = cfgOut[38:36]; // @[PE.scala 113:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 70:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_1_io_config = cfgOut[41:39]; // @[PE.scala 113:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 70:23]
  assign Muxn_io_config = cfgOut[44:42]; // @[PE.scala 121:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 62:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 62:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 62:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 62:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign Muxn_1_io_config = cfgOut[47:45]; // @[PE.scala 121:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 62:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 62:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 62:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 62:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 90:17]
  assign cfg_io_cfg_addr = io_cfg_addr[0]; // @[PE.scala 91:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 92:19]
endmodule
module GPE_9(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [3:0] alu_io_config; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 50:19]
  wire [31:0] alu_io_out; // @[PE.scala 50:19]
  wire  rf_clock; // @[PE.scala 51:18]
  wire  rf_reset; // @[PE.scala 51:18]
  wire  rf_io_en; // @[PE.scala 51:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 51:18]
  wire  DelayPipe_clock; // @[PE.scala 52:54]
  wire  DelayPipe_reset; // @[PE.scala 52:54]
  wire  DelayPipe_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 52:54]
  wire  DelayPipe_1_clock; // @[PE.scala 52:54]
  wire  DelayPipe_1_reset; // @[PE.scala 52:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 52:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 55:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 55:49]
  wire  cfg_clock; // @[PE.scala 89:19]
  wire  cfg_reset; // @[PE.scala 89:19]
  wire  cfg_io_cfg_en; // @[PE.scala 89:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 89:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 89:19]
  wire [47:0] cfg_io_out_0; // @[PE.scala 89:19]
  wire  _T_1 = 10'h2f == io_cfg_addr[11:2]; // @[PE.scala 90:48]
  wire [47:0] cfgOut = cfg_io_out_0; // @[PE.scala 96:20 PE.scala 97:10]
  ALU alu ( // @[PE.scala 50:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 51:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 52:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 52:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_16 Muxn ( // @[PE.scala 55:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_16 Muxn_1 ( // @[PE.scala 55:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_16 cfg ( // @[PE.scala 89:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 77:13]
  assign alu_io_config = cfgOut[35:32]; // @[PE.scala 100:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 71:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 71:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 75:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 76:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_io_config = cfgOut[38:36]; // @[PE.scala 113:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 70:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_1_io_config = cfgOut[41:39]; // @[PE.scala 113:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 70:23]
  assign Muxn_io_config = cfgOut[44:42]; // @[PE.scala 121:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 62:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 62:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 62:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 62:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign Muxn_1_io_config = cfgOut[47:45]; // @[PE.scala 121:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 62:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 62:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 62:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 62:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 90:17]
  assign cfg_io_cfg_addr = io_cfg_addr[0]; // @[PE.scala 91:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 92:19]
endmodule
module GPE_10(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [3:0] alu_io_config; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 50:19]
  wire [31:0] alu_io_out; // @[PE.scala 50:19]
  wire  rf_clock; // @[PE.scala 51:18]
  wire  rf_reset; // @[PE.scala 51:18]
  wire  rf_io_en; // @[PE.scala 51:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 51:18]
  wire  DelayPipe_clock; // @[PE.scala 52:54]
  wire  DelayPipe_reset; // @[PE.scala 52:54]
  wire  DelayPipe_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 52:54]
  wire  DelayPipe_1_clock; // @[PE.scala 52:54]
  wire  DelayPipe_1_reset; // @[PE.scala 52:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 52:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 55:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 55:49]
  wire  cfg_clock; // @[PE.scala 89:19]
  wire  cfg_reset; // @[PE.scala 89:19]
  wire  cfg_io_cfg_en; // @[PE.scala 89:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 89:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 89:19]
  wire [47:0] cfg_io_out_0; // @[PE.scala 89:19]
  wire  _T_1 = 10'h30 == io_cfg_addr[11:2]; // @[PE.scala 90:48]
  wire [47:0] cfgOut = cfg_io_out_0; // @[PE.scala 96:20 PE.scala 97:10]
  ALU alu ( // @[PE.scala 50:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 51:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 52:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 52:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_16 Muxn ( // @[PE.scala 55:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_16 Muxn_1 ( // @[PE.scala 55:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_16 cfg ( // @[PE.scala 89:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 77:13]
  assign alu_io_config = cfgOut[35:32]; // @[PE.scala 100:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 71:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 71:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 75:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 76:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_io_config = cfgOut[38:36]; // @[PE.scala 113:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 70:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_1_io_config = cfgOut[41:39]; // @[PE.scala 113:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 70:23]
  assign Muxn_io_config = cfgOut[44:42]; // @[PE.scala 121:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 62:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 62:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 62:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 62:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign Muxn_1_io_config = cfgOut[47:45]; // @[PE.scala 121:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 62:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 62:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 62:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 62:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 90:17]
  assign cfg_io_cfg_addr = io_cfg_addr[0]; // @[PE.scala 91:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 92:19]
endmodule
module GPE_11(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [3:0] alu_io_config; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 50:19]
  wire [31:0] alu_io_out; // @[PE.scala 50:19]
  wire  rf_clock; // @[PE.scala 51:18]
  wire  rf_reset; // @[PE.scala 51:18]
  wire  rf_io_en; // @[PE.scala 51:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 51:18]
  wire  DelayPipe_clock; // @[PE.scala 52:54]
  wire  DelayPipe_reset; // @[PE.scala 52:54]
  wire  DelayPipe_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 52:54]
  wire  DelayPipe_1_clock; // @[PE.scala 52:54]
  wire  DelayPipe_1_reset; // @[PE.scala 52:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 52:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 55:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 55:49]
  wire  cfg_clock; // @[PE.scala 89:19]
  wire  cfg_reset; // @[PE.scala 89:19]
  wire  cfg_io_cfg_en; // @[PE.scala 89:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 89:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 89:19]
  wire [47:0] cfg_io_out_0; // @[PE.scala 89:19]
  wire  _T_1 = 10'h31 == io_cfg_addr[11:2]; // @[PE.scala 90:48]
  wire [47:0] cfgOut = cfg_io_out_0; // @[PE.scala 96:20 PE.scala 97:10]
  ALU alu ( // @[PE.scala 50:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 51:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 52:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 52:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_16 Muxn ( // @[PE.scala 55:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_16 Muxn_1 ( // @[PE.scala 55:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_16 cfg ( // @[PE.scala 89:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 77:13]
  assign alu_io_config = cfgOut[35:32]; // @[PE.scala 100:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 71:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 71:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 75:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 76:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_io_config = cfgOut[38:36]; // @[PE.scala 113:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 70:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_1_io_config = cfgOut[41:39]; // @[PE.scala 113:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 70:23]
  assign Muxn_io_config = cfgOut[44:42]; // @[PE.scala 121:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 62:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 62:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 62:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 62:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign Muxn_1_io_config = cfgOut[47:45]; // @[PE.scala 121:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 62:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 62:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 62:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 62:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 90:17]
  assign cfg_io_cfg_addr = io_cfg_addr[0]; // @[PE.scala 91:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 92:19]
endmodule
module GPE_12(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [3:0] alu_io_config; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 50:19]
  wire [31:0] alu_io_out; // @[PE.scala 50:19]
  wire  rf_clock; // @[PE.scala 51:18]
  wire  rf_reset; // @[PE.scala 51:18]
  wire  rf_io_en; // @[PE.scala 51:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 51:18]
  wire  DelayPipe_clock; // @[PE.scala 52:54]
  wire  DelayPipe_reset; // @[PE.scala 52:54]
  wire  DelayPipe_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 52:54]
  wire  DelayPipe_1_clock; // @[PE.scala 52:54]
  wire  DelayPipe_1_reset; // @[PE.scala 52:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 52:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 55:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 55:49]
  wire  cfg_clock; // @[PE.scala 89:19]
  wire  cfg_reset; // @[PE.scala 89:19]
  wire  cfg_io_cfg_en; // @[PE.scala 89:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 89:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 89:19]
  wire [47:0] cfg_io_out_0; // @[PE.scala 89:19]
  wire  _T_1 = 10'h32 == io_cfg_addr[11:2]; // @[PE.scala 90:48]
  wire [47:0] cfgOut = cfg_io_out_0; // @[PE.scala 96:20 PE.scala 97:10]
  ALU alu ( // @[PE.scala 50:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 51:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 52:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 52:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_16 Muxn ( // @[PE.scala 55:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_16 Muxn_1 ( // @[PE.scala 55:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_16 cfg ( // @[PE.scala 89:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 77:13]
  assign alu_io_config = cfgOut[35:32]; // @[PE.scala 100:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 71:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 71:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 75:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 76:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_io_config = cfgOut[38:36]; // @[PE.scala 113:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 70:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_1_io_config = cfgOut[41:39]; // @[PE.scala 113:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 70:23]
  assign Muxn_io_config = cfgOut[44:42]; // @[PE.scala 121:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 62:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 62:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 62:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 62:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign Muxn_1_io_config = cfgOut[47:45]; // @[PE.scala 121:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 62:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 62:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 62:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 62:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 90:17]
  assign cfg_io_cfg_addr = io_cfg_addr[0]; // @[PE.scala 91:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 92:19]
endmodule
module GPE_13(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [3:0] alu_io_config; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 50:19]
  wire [31:0] alu_io_out; // @[PE.scala 50:19]
  wire  rf_clock; // @[PE.scala 51:18]
  wire  rf_reset; // @[PE.scala 51:18]
  wire  rf_io_en; // @[PE.scala 51:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 51:18]
  wire  DelayPipe_clock; // @[PE.scala 52:54]
  wire  DelayPipe_reset; // @[PE.scala 52:54]
  wire  DelayPipe_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 52:54]
  wire  DelayPipe_1_clock; // @[PE.scala 52:54]
  wire  DelayPipe_1_reset; // @[PE.scala 52:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 52:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 55:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 55:49]
  wire  cfg_clock; // @[PE.scala 89:19]
  wire  cfg_reset; // @[PE.scala 89:19]
  wire  cfg_io_cfg_en; // @[PE.scala 89:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 89:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 89:19]
  wire [47:0] cfg_io_out_0; // @[PE.scala 89:19]
  wire  _T_1 = 10'h33 == io_cfg_addr[11:2]; // @[PE.scala 90:48]
  wire [47:0] cfgOut = cfg_io_out_0; // @[PE.scala 96:20 PE.scala 97:10]
  ALU alu ( // @[PE.scala 50:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 51:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 52:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 52:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_16 Muxn ( // @[PE.scala 55:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_16 Muxn_1 ( // @[PE.scala 55:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_16 cfg ( // @[PE.scala 89:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 77:13]
  assign alu_io_config = cfgOut[35:32]; // @[PE.scala 100:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 71:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 71:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 75:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 76:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_io_config = cfgOut[38:36]; // @[PE.scala 113:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 70:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_1_io_config = cfgOut[41:39]; // @[PE.scala 113:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 70:23]
  assign Muxn_io_config = cfgOut[44:42]; // @[PE.scala 121:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 62:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 62:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 62:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 62:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign Muxn_1_io_config = cfgOut[47:45]; // @[PE.scala 121:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 62:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 62:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 62:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 62:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 90:17]
  assign cfg_io_cfg_addr = io_cfg_addr[0]; // @[PE.scala 91:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 92:19]
endmodule
module GPE_14(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [3:0] alu_io_config; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 50:19]
  wire [31:0] alu_io_out; // @[PE.scala 50:19]
  wire  rf_clock; // @[PE.scala 51:18]
  wire  rf_reset; // @[PE.scala 51:18]
  wire  rf_io_en; // @[PE.scala 51:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 51:18]
  wire  DelayPipe_clock; // @[PE.scala 52:54]
  wire  DelayPipe_reset; // @[PE.scala 52:54]
  wire  DelayPipe_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 52:54]
  wire  DelayPipe_1_clock; // @[PE.scala 52:54]
  wire  DelayPipe_1_reset; // @[PE.scala 52:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 52:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 55:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 55:49]
  wire  cfg_clock; // @[PE.scala 89:19]
  wire  cfg_reset; // @[PE.scala 89:19]
  wire  cfg_io_cfg_en; // @[PE.scala 89:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 89:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 89:19]
  wire [47:0] cfg_io_out_0; // @[PE.scala 89:19]
  wire  _T_1 = 10'h34 == io_cfg_addr[11:2]; // @[PE.scala 90:48]
  wire [47:0] cfgOut = cfg_io_out_0; // @[PE.scala 96:20 PE.scala 97:10]
  ALU alu ( // @[PE.scala 50:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 51:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 52:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 52:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_16 Muxn ( // @[PE.scala 55:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_16 Muxn_1 ( // @[PE.scala 55:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_16 cfg ( // @[PE.scala 89:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 77:13]
  assign alu_io_config = cfgOut[35:32]; // @[PE.scala 100:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 71:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 71:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 75:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 76:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_io_config = cfgOut[38:36]; // @[PE.scala 113:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 70:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_1_io_config = cfgOut[41:39]; // @[PE.scala 113:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 70:23]
  assign Muxn_io_config = cfgOut[44:42]; // @[PE.scala 121:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 62:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 62:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 62:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 62:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign Muxn_1_io_config = cfgOut[47:45]; // @[PE.scala 121:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 62:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 62:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 62:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 62:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 90:17]
  assign cfg_io_cfg_addr = io_cfg_addr[0]; // @[PE.scala 91:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 92:19]
endmodule
module GPE_15(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [3:0] alu_io_config; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 50:19]
  wire [31:0] alu_io_out; // @[PE.scala 50:19]
  wire  rf_clock; // @[PE.scala 51:18]
  wire  rf_reset; // @[PE.scala 51:18]
  wire  rf_io_en; // @[PE.scala 51:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 51:18]
  wire  DelayPipe_clock; // @[PE.scala 52:54]
  wire  DelayPipe_reset; // @[PE.scala 52:54]
  wire  DelayPipe_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 52:54]
  wire  DelayPipe_1_clock; // @[PE.scala 52:54]
  wire  DelayPipe_1_reset; // @[PE.scala 52:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 52:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 55:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 55:49]
  wire  cfg_clock; // @[PE.scala 89:19]
  wire  cfg_reset; // @[PE.scala 89:19]
  wire  cfg_io_cfg_en; // @[PE.scala 89:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 89:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 89:19]
  wire [47:0] cfg_io_out_0; // @[PE.scala 89:19]
  wire  _T_1 = 10'h35 == io_cfg_addr[11:2]; // @[PE.scala 90:48]
  wire [47:0] cfgOut = cfg_io_out_0; // @[PE.scala 96:20 PE.scala 97:10]
  ALU alu ( // @[PE.scala 50:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 51:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 52:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 52:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_16 Muxn ( // @[PE.scala 55:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_16 Muxn_1 ( // @[PE.scala 55:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_16 cfg ( // @[PE.scala 89:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 77:13]
  assign alu_io_config = cfgOut[35:32]; // @[PE.scala 100:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 71:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 71:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 75:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 76:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_io_config = cfgOut[38:36]; // @[PE.scala 113:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 70:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_1_io_config = cfgOut[41:39]; // @[PE.scala 113:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 70:23]
  assign Muxn_io_config = cfgOut[44:42]; // @[PE.scala 121:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 62:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 62:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 62:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 62:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign Muxn_1_io_config = cfgOut[47:45]; // @[PE.scala 121:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 62:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 62:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 62:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 62:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 90:17]
  assign cfg_io_cfg_addr = io_cfg_addr[0]; // @[PE.scala 91:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 92:19]
endmodule
module GPE_16(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [3:0] alu_io_config; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 50:19]
  wire [31:0] alu_io_out; // @[PE.scala 50:19]
  wire  rf_clock; // @[PE.scala 51:18]
  wire  rf_reset; // @[PE.scala 51:18]
  wire  rf_io_en; // @[PE.scala 51:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 51:18]
  wire  DelayPipe_clock; // @[PE.scala 52:54]
  wire  DelayPipe_reset; // @[PE.scala 52:54]
  wire  DelayPipe_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 52:54]
  wire  DelayPipe_1_clock; // @[PE.scala 52:54]
  wire  DelayPipe_1_reset; // @[PE.scala 52:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 52:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 55:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 55:49]
  wire  cfg_clock; // @[PE.scala 89:19]
  wire  cfg_reset; // @[PE.scala 89:19]
  wire  cfg_io_cfg_en; // @[PE.scala 89:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 89:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 89:19]
  wire [47:0] cfg_io_out_0; // @[PE.scala 89:19]
  wire  _T_1 = 10'h40 == io_cfg_addr[11:2]; // @[PE.scala 90:48]
  wire [47:0] cfgOut = cfg_io_out_0; // @[PE.scala 96:20 PE.scala 97:10]
  ALU alu ( // @[PE.scala 50:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 51:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 52:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 52:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_16 Muxn ( // @[PE.scala 55:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_16 Muxn_1 ( // @[PE.scala 55:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_16 cfg ( // @[PE.scala 89:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 77:13]
  assign alu_io_config = cfgOut[35:32]; // @[PE.scala 100:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 71:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 71:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 75:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 76:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_io_config = cfgOut[38:36]; // @[PE.scala 113:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 70:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_1_io_config = cfgOut[41:39]; // @[PE.scala 113:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 70:23]
  assign Muxn_io_config = cfgOut[44:42]; // @[PE.scala 121:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 62:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 62:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 62:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 62:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign Muxn_1_io_config = cfgOut[47:45]; // @[PE.scala 121:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 62:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 62:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 62:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 62:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 90:17]
  assign cfg_io_cfg_addr = io_cfg_addr[0]; // @[PE.scala 91:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 92:19]
endmodule
module GPE_17(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [3:0] alu_io_config; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 50:19]
  wire [31:0] alu_io_out; // @[PE.scala 50:19]
  wire  rf_clock; // @[PE.scala 51:18]
  wire  rf_reset; // @[PE.scala 51:18]
  wire  rf_io_en; // @[PE.scala 51:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 51:18]
  wire  DelayPipe_clock; // @[PE.scala 52:54]
  wire  DelayPipe_reset; // @[PE.scala 52:54]
  wire  DelayPipe_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 52:54]
  wire  DelayPipe_1_clock; // @[PE.scala 52:54]
  wire  DelayPipe_1_reset; // @[PE.scala 52:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 52:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 55:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 55:49]
  wire  cfg_clock; // @[PE.scala 89:19]
  wire  cfg_reset; // @[PE.scala 89:19]
  wire  cfg_io_cfg_en; // @[PE.scala 89:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 89:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 89:19]
  wire [47:0] cfg_io_out_0; // @[PE.scala 89:19]
  wire  _T_1 = 10'h41 == io_cfg_addr[11:2]; // @[PE.scala 90:48]
  wire [47:0] cfgOut = cfg_io_out_0; // @[PE.scala 96:20 PE.scala 97:10]
  ALU alu ( // @[PE.scala 50:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 51:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 52:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 52:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_16 Muxn ( // @[PE.scala 55:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_16 Muxn_1 ( // @[PE.scala 55:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_16 cfg ( // @[PE.scala 89:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 77:13]
  assign alu_io_config = cfgOut[35:32]; // @[PE.scala 100:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 71:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 71:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 75:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 76:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_io_config = cfgOut[38:36]; // @[PE.scala 113:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 70:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_1_io_config = cfgOut[41:39]; // @[PE.scala 113:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 70:23]
  assign Muxn_io_config = cfgOut[44:42]; // @[PE.scala 121:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 62:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 62:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 62:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 62:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign Muxn_1_io_config = cfgOut[47:45]; // @[PE.scala 121:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 62:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 62:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 62:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 62:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 90:17]
  assign cfg_io_cfg_addr = io_cfg_addr[0]; // @[PE.scala 91:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 92:19]
endmodule
module GPE_18(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [3:0] alu_io_config; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 50:19]
  wire [31:0] alu_io_out; // @[PE.scala 50:19]
  wire  rf_clock; // @[PE.scala 51:18]
  wire  rf_reset; // @[PE.scala 51:18]
  wire  rf_io_en; // @[PE.scala 51:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 51:18]
  wire  DelayPipe_clock; // @[PE.scala 52:54]
  wire  DelayPipe_reset; // @[PE.scala 52:54]
  wire  DelayPipe_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 52:54]
  wire  DelayPipe_1_clock; // @[PE.scala 52:54]
  wire  DelayPipe_1_reset; // @[PE.scala 52:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 52:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 55:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 55:49]
  wire  cfg_clock; // @[PE.scala 89:19]
  wire  cfg_reset; // @[PE.scala 89:19]
  wire  cfg_io_cfg_en; // @[PE.scala 89:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 89:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 89:19]
  wire [47:0] cfg_io_out_0; // @[PE.scala 89:19]
  wire  _T_1 = 10'h42 == io_cfg_addr[11:2]; // @[PE.scala 90:48]
  wire [47:0] cfgOut = cfg_io_out_0; // @[PE.scala 96:20 PE.scala 97:10]
  ALU alu ( // @[PE.scala 50:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 51:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 52:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 52:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_16 Muxn ( // @[PE.scala 55:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_16 Muxn_1 ( // @[PE.scala 55:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_16 cfg ( // @[PE.scala 89:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 77:13]
  assign alu_io_config = cfgOut[35:32]; // @[PE.scala 100:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 71:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 71:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 75:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 76:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_io_config = cfgOut[38:36]; // @[PE.scala 113:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 70:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_1_io_config = cfgOut[41:39]; // @[PE.scala 113:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 70:23]
  assign Muxn_io_config = cfgOut[44:42]; // @[PE.scala 121:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 62:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 62:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 62:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 62:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign Muxn_1_io_config = cfgOut[47:45]; // @[PE.scala 121:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 62:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 62:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 62:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 62:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 90:17]
  assign cfg_io_cfg_addr = io_cfg_addr[0]; // @[PE.scala 91:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 92:19]
endmodule
module GPE_19(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [3:0] alu_io_config; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 50:19]
  wire [31:0] alu_io_out; // @[PE.scala 50:19]
  wire  rf_clock; // @[PE.scala 51:18]
  wire  rf_reset; // @[PE.scala 51:18]
  wire  rf_io_en; // @[PE.scala 51:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 51:18]
  wire  DelayPipe_clock; // @[PE.scala 52:54]
  wire  DelayPipe_reset; // @[PE.scala 52:54]
  wire  DelayPipe_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 52:54]
  wire  DelayPipe_1_clock; // @[PE.scala 52:54]
  wire  DelayPipe_1_reset; // @[PE.scala 52:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 52:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 55:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 55:49]
  wire  cfg_clock; // @[PE.scala 89:19]
  wire  cfg_reset; // @[PE.scala 89:19]
  wire  cfg_io_cfg_en; // @[PE.scala 89:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 89:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 89:19]
  wire [47:0] cfg_io_out_0; // @[PE.scala 89:19]
  wire  _T_1 = 10'h43 == io_cfg_addr[11:2]; // @[PE.scala 90:48]
  wire [47:0] cfgOut = cfg_io_out_0; // @[PE.scala 96:20 PE.scala 97:10]
  ALU alu ( // @[PE.scala 50:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 51:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 52:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 52:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_16 Muxn ( // @[PE.scala 55:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_16 Muxn_1 ( // @[PE.scala 55:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_16 cfg ( // @[PE.scala 89:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 77:13]
  assign alu_io_config = cfgOut[35:32]; // @[PE.scala 100:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 71:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 71:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 75:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 76:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_io_config = cfgOut[38:36]; // @[PE.scala 113:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 70:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_1_io_config = cfgOut[41:39]; // @[PE.scala 113:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 70:23]
  assign Muxn_io_config = cfgOut[44:42]; // @[PE.scala 121:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 62:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 62:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 62:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 62:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign Muxn_1_io_config = cfgOut[47:45]; // @[PE.scala 121:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 62:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 62:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 62:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 62:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 90:17]
  assign cfg_io_cfg_addr = io_cfg_addr[0]; // @[PE.scala 91:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 92:19]
endmodule
module GPE_20(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [3:0] alu_io_config; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 50:19]
  wire [31:0] alu_io_out; // @[PE.scala 50:19]
  wire  rf_clock; // @[PE.scala 51:18]
  wire  rf_reset; // @[PE.scala 51:18]
  wire  rf_io_en; // @[PE.scala 51:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 51:18]
  wire  DelayPipe_clock; // @[PE.scala 52:54]
  wire  DelayPipe_reset; // @[PE.scala 52:54]
  wire  DelayPipe_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 52:54]
  wire  DelayPipe_1_clock; // @[PE.scala 52:54]
  wire  DelayPipe_1_reset; // @[PE.scala 52:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 52:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 55:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 55:49]
  wire  cfg_clock; // @[PE.scala 89:19]
  wire  cfg_reset; // @[PE.scala 89:19]
  wire  cfg_io_cfg_en; // @[PE.scala 89:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 89:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 89:19]
  wire [47:0] cfg_io_out_0; // @[PE.scala 89:19]
  wire  _T_1 = 10'h44 == io_cfg_addr[11:2]; // @[PE.scala 90:48]
  wire [47:0] cfgOut = cfg_io_out_0; // @[PE.scala 96:20 PE.scala 97:10]
  ALU alu ( // @[PE.scala 50:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 51:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 52:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 52:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_16 Muxn ( // @[PE.scala 55:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_16 Muxn_1 ( // @[PE.scala 55:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_16 cfg ( // @[PE.scala 89:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 77:13]
  assign alu_io_config = cfgOut[35:32]; // @[PE.scala 100:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 71:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 71:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 75:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 76:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_io_config = cfgOut[38:36]; // @[PE.scala 113:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 70:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_1_io_config = cfgOut[41:39]; // @[PE.scala 113:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 70:23]
  assign Muxn_io_config = cfgOut[44:42]; // @[PE.scala 121:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 62:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 62:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 62:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 62:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign Muxn_1_io_config = cfgOut[47:45]; // @[PE.scala 121:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 62:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 62:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 62:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 62:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 90:17]
  assign cfg_io_cfg_addr = io_cfg_addr[0]; // @[PE.scala 91:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 92:19]
endmodule
module GPE_21(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [3:0] alu_io_config; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 50:19]
  wire [31:0] alu_io_out; // @[PE.scala 50:19]
  wire  rf_clock; // @[PE.scala 51:18]
  wire  rf_reset; // @[PE.scala 51:18]
  wire  rf_io_en; // @[PE.scala 51:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 51:18]
  wire  DelayPipe_clock; // @[PE.scala 52:54]
  wire  DelayPipe_reset; // @[PE.scala 52:54]
  wire  DelayPipe_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 52:54]
  wire  DelayPipe_1_clock; // @[PE.scala 52:54]
  wire  DelayPipe_1_reset; // @[PE.scala 52:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 52:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 55:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 55:49]
  wire  cfg_clock; // @[PE.scala 89:19]
  wire  cfg_reset; // @[PE.scala 89:19]
  wire  cfg_io_cfg_en; // @[PE.scala 89:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 89:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 89:19]
  wire [47:0] cfg_io_out_0; // @[PE.scala 89:19]
  wire  _T_1 = 10'h45 == io_cfg_addr[11:2]; // @[PE.scala 90:48]
  wire [47:0] cfgOut = cfg_io_out_0; // @[PE.scala 96:20 PE.scala 97:10]
  ALU alu ( // @[PE.scala 50:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 51:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 52:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 52:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_16 Muxn ( // @[PE.scala 55:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_16 Muxn_1 ( // @[PE.scala 55:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_16 cfg ( // @[PE.scala 89:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 77:13]
  assign alu_io_config = cfgOut[35:32]; // @[PE.scala 100:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 71:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 71:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 75:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 76:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_io_config = cfgOut[38:36]; // @[PE.scala 113:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 70:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_1_io_config = cfgOut[41:39]; // @[PE.scala 113:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 70:23]
  assign Muxn_io_config = cfgOut[44:42]; // @[PE.scala 121:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 62:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 62:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 62:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 62:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign Muxn_1_io_config = cfgOut[47:45]; // @[PE.scala 121:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 62:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 62:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 62:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 62:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 90:17]
  assign cfg_io_cfg_addr = io_cfg_addr[0]; // @[PE.scala 91:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 92:19]
endmodule
module GPE_22(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [3:0] alu_io_config; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 50:19]
  wire [31:0] alu_io_out; // @[PE.scala 50:19]
  wire  rf_clock; // @[PE.scala 51:18]
  wire  rf_reset; // @[PE.scala 51:18]
  wire  rf_io_en; // @[PE.scala 51:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 51:18]
  wire  DelayPipe_clock; // @[PE.scala 52:54]
  wire  DelayPipe_reset; // @[PE.scala 52:54]
  wire  DelayPipe_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 52:54]
  wire  DelayPipe_1_clock; // @[PE.scala 52:54]
  wire  DelayPipe_1_reset; // @[PE.scala 52:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 52:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 55:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 55:49]
  wire  cfg_clock; // @[PE.scala 89:19]
  wire  cfg_reset; // @[PE.scala 89:19]
  wire  cfg_io_cfg_en; // @[PE.scala 89:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 89:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 89:19]
  wire [47:0] cfg_io_out_0; // @[PE.scala 89:19]
  wire  _T_1 = 10'h46 == io_cfg_addr[11:2]; // @[PE.scala 90:48]
  wire [47:0] cfgOut = cfg_io_out_0; // @[PE.scala 96:20 PE.scala 97:10]
  ALU alu ( // @[PE.scala 50:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 51:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 52:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 52:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_16 Muxn ( // @[PE.scala 55:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_16 Muxn_1 ( // @[PE.scala 55:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_16 cfg ( // @[PE.scala 89:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 77:13]
  assign alu_io_config = cfgOut[35:32]; // @[PE.scala 100:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 71:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 71:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 75:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 76:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_io_config = cfgOut[38:36]; // @[PE.scala 113:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 70:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_1_io_config = cfgOut[41:39]; // @[PE.scala 113:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 70:23]
  assign Muxn_io_config = cfgOut[44:42]; // @[PE.scala 121:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 62:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 62:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 62:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 62:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign Muxn_1_io_config = cfgOut[47:45]; // @[PE.scala 121:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 62:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 62:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 62:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 62:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 90:17]
  assign cfg_io_cfg_addr = io_cfg_addr[0]; // @[PE.scala 91:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 92:19]
endmodule
module GPE_23(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [3:0] alu_io_config; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 50:19]
  wire [31:0] alu_io_out; // @[PE.scala 50:19]
  wire  rf_clock; // @[PE.scala 51:18]
  wire  rf_reset; // @[PE.scala 51:18]
  wire  rf_io_en; // @[PE.scala 51:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 51:18]
  wire  DelayPipe_clock; // @[PE.scala 52:54]
  wire  DelayPipe_reset; // @[PE.scala 52:54]
  wire  DelayPipe_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 52:54]
  wire  DelayPipe_1_clock; // @[PE.scala 52:54]
  wire  DelayPipe_1_reset; // @[PE.scala 52:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 52:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 55:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 55:49]
  wire  cfg_clock; // @[PE.scala 89:19]
  wire  cfg_reset; // @[PE.scala 89:19]
  wire  cfg_io_cfg_en; // @[PE.scala 89:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 89:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 89:19]
  wire [47:0] cfg_io_out_0; // @[PE.scala 89:19]
  wire  _T_1 = 10'h47 == io_cfg_addr[11:2]; // @[PE.scala 90:48]
  wire [47:0] cfgOut = cfg_io_out_0; // @[PE.scala 96:20 PE.scala 97:10]
  ALU alu ( // @[PE.scala 50:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 51:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 52:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 52:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_16 Muxn ( // @[PE.scala 55:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_16 Muxn_1 ( // @[PE.scala 55:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_16 cfg ( // @[PE.scala 89:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 77:13]
  assign alu_io_config = cfgOut[35:32]; // @[PE.scala 100:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 71:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 71:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 75:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 76:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_io_config = cfgOut[38:36]; // @[PE.scala 113:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 70:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_1_io_config = cfgOut[41:39]; // @[PE.scala 113:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 70:23]
  assign Muxn_io_config = cfgOut[44:42]; // @[PE.scala 121:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 62:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 62:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 62:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 62:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign Muxn_1_io_config = cfgOut[47:45]; // @[PE.scala 121:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 62:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 62:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 62:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 62:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 90:17]
  assign cfg_io_cfg_addr = io_cfg_addr[0]; // @[PE.scala 91:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 92:19]
endmodule
module GPE_24(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [3:0] alu_io_config; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 50:19]
  wire [31:0] alu_io_out; // @[PE.scala 50:19]
  wire  rf_clock; // @[PE.scala 51:18]
  wire  rf_reset; // @[PE.scala 51:18]
  wire  rf_io_en; // @[PE.scala 51:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 51:18]
  wire  DelayPipe_clock; // @[PE.scala 52:54]
  wire  DelayPipe_reset; // @[PE.scala 52:54]
  wire  DelayPipe_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 52:54]
  wire  DelayPipe_1_clock; // @[PE.scala 52:54]
  wire  DelayPipe_1_reset; // @[PE.scala 52:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 52:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 55:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 55:49]
  wire  cfg_clock; // @[PE.scala 89:19]
  wire  cfg_reset; // @[PE.scala 89:19]
  wire  cfg_io_cfg_en; // @[PE.scala 89:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 89:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 89:19]
  wire [47:0] cfg_io_out_0; // @[PE.scala 89:19]
  wire  _T_1 = 10'h52 == io_cfg_addr[11:2]; // @[PE.scala 90:48]
  wire [47:0] cfgOut = cfg_io_out_0; // @[PE.scala 96:20 PE.scala 97:10]
  ALU alu ( // @[PE.scala 50:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 51:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 52:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 52:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_16 Muxn ( // @[PE.scala 55:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_16 Muxn_1 ( // @[PE.scala 55:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_16 cfg ( // @[PE.scala 89:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 77:13]
  assign alu_io_config = cfgOut[35:32]; // @[PE.scala 100:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 71:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 71:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 75:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 76:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_io_config = cfgOut[38:36]; // @[PE.scala 113:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 70:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_1_io_config = cfgOut[41:39]; // @[PE.scala 113:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 70:23]
  assign Muxn_io_config = cfgOut[44:42]; // @[PE.scala 121:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 62:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 62:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 62:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 62:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign Muxn_1_io_config = cfgOut[47:45]; // @[PE.scala 121:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 62:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 62:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 62:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 62:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 90:17]
  assign cfg_io_cfg_addr = io_cfg_addr[0]; // @[PE.scala 91:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 92:19]
endmodule
module GPE_25(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [3:0] alu_io_config; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 50:19]
  wire [31:0] alu_io_out; // @[PE.scala 50:19]
  wire  rf_clock; // @[PE.scala 51:18]
  wire  rf_reset; // @[PE.scala 51:18]
  wire  rf_io_en; // @[PE.scala 51:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 51:18]
  wire  DelayPipe_clock; // @[PE.scala 52:54]
  wire  DelayPipe_reset; // @[PE.scala 52:54]
  wire  DelayPipe_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 52:54]
  wire  DelayPipe_1_clock; // @[PE.scala 52:54]
  wire  DelayPipe_1_reset; // @[PE.scala 52:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 52:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 55:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 55:49]
  wire  cfg_clock; // @[PE.scala 89:19]
  wire  cfg_reset; // @[PE.scala 89:19]
  wire  cfg_io_cfg_en; // @[PE.scala 89:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 89:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 89:19]
  wire [47:0] cfg_io_out_0; // @[PE.scala 89:19]
  wire  _T_1 = 10'h53 == io_cfg_addr[11:2]; // @[PE.scala 90:48]
  wire [47:0] cfgOut = cfg_io_out_0; // @[PE.scala 96:20 PE.scala 97:10]
  ALU alu ( // @[PE.scala 50:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 51:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 52:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 52:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_16 Muxn ( // @[PE.scala 55:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_16 Muxn_1 ( // @[PE.scala 55:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_16 cfg ( // @[PE.scala 89:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 77:13]
  assign alu_io_config = cfgOut[35:32]; // @[PE.scala 100:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 71:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 71:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 75:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 76:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_io_config = cfgOut[38:36]; // @[PE.scala 113:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 70:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_1_io_config = cfgOut[41:39]; // @[PE.scala 113:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 70:23]
  assign Muxn_io_config = cfgOut[44:42]; // @[PE.scala 121:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 62:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 62:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 62:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 62:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign Muxn_1_io_config = cfgOut[47:45]; // @[PE.scala 121:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 62:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 62:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 62:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 62:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 90:17]
  assign cfg_io_cfg_addr = io_cfg_addr[0]; // @[PE.scala 91:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 92:19]
endmodule
module GPE_26(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [3:0] alu_io_config; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 50:19]
  wire [31:0] alu_io_out; // @[PE.scala 50:19]
  wire  rf_clock; // @[PE.scala 51:18]
  wire  rf_reset; // @[PE.scala 51:18]
  wire  rf_io_en; // @[PE.scala 51:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 51:18]
  wire  DelayPipe_clock; // @[PE.scala 52:54]
  wire  DelayPipe_reset; // @[PE.scala 52:54]
  wire  DelayPipe_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 52:54]
  wire  DelayPipe_1_clock; // @[PE.scala 52:54]
  wire  DelayPipe_1_reset; // @[PE.scala 52:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 52:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 55:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 55:49]
  wire  cfg_clock; // @[PE.scala 89:19]
  wire  cfg_reset; // @[PE.scala 89:19]
  wire  cfg_io_cfg_en; // @[PE.scala 89:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 89:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 89:19]
  wire [47:0] cfg_io_out_0; // @[PE.scala 89:19]
  wire  _T_1 = 10'h54 == io_cfg_addr[11:2]; // @[PE.scala 90:48]
  wire [47:0] cfgOut = cfg_io_out_0; // @[PE.scala 96:20 PE.scala 97:10]
  ALU alu ( // @[PE.scala 50:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 51:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 52:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 52:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_16 Muxn ( // @[PE.scala 55:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_16 Muxn_1 ( // @[PE.scala 55:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_16 cfg ( // @[PE.scala 89:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 77:13]
  assign alu_io_config = cfgOut[35:32]; // @[PE.scala 100:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 71:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 71:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 75:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 76:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_io_config = cfgOut[38:36]; // @[PE.scala 113:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 70:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_1_io_config = cfgOut[41:39]; // @[PE.scala 113:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 70:23]
  assign Muxn_io_config = cfgOut[44:42]; // @[PE.scala 121:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 62:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 62:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 62:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 62:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign Muxn_1_io_config = cfgOut[47:45]; // @[PE.scala 121:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 62:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 62:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 62:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 62:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 90:17]
  assign cfg_io_cfg_addr = io_cfg_addr[0]; // @[PE.scala 91:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 92:19]
endmodule
module GPE_27(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [3:0] alu_io_config; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 50:19]
  wire [31:0] alu_io_out; // @[PE.scala 50:19]
  wire  rf_clock; // @[PE.scala 51:18]
  wire  rf_reset; // @[PE.scala 51:18]
  wire  rf_io_en; // @[PE.scala 51:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 51:18]
  wire  DelayPipe_clock; // @[PE.scala 52:54]
  wire  DelayPipe_reset; // @[PE.scala 52:54]
  wire  DelayPipe_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 52:54]
  wire  DelayPipe_1_clock; // @[PE.scala 52:54]
  wire  DelayPipe_1_reset; // @[PE.scala 52:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 52:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 55:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 55:49]
  wire  cfg_clock; // @[PE.scala 89:19]
  wire  cfg_reset; // @[PE.scala 89:19]
  wire  cfg_io_cfg_en; // @[PE.scala 89:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 89:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 89:19]
  wire [47:0] cfg_io_out_0; // @[PE.scala 89:19]
  wire  _T_1 = 10'h55 == io_cfg_addr[11:2]; // @[PE.scala 90:48]
  wire [47:0] cfgOut = cfg_io_out_0; // @[PE.scala 96:20 PE.scala 97:10]
  ALU alu ( // @[PE.scala 50:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 51:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 52:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 52:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_16 Muxn ( // @[PE.scala 55:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_16 Muxn_1 ( // @[PE.scala 55:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_16 cfg ( // @[PE.scala 89:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 77:13]
  assign alu_io_config = cfgOut[35:32]; // @[PE.scala 100:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 71:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 71:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 75:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 76:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_io_config = cfgOut[38:36]; // @[PE.scala 113:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 70:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_1_io_config = cfgOut[41:39]; // @[PE.scala 113:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 70:23]
  assign Muxn_io_config = cfgOut[44:42]; // @[PE.scala 121:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 62:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 62:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 62:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 62:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign Muxn_1_io_config = cfgOut[47:45]; // @[PE.scala 121:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 62:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 62:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 62:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 62:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 90:17]
  assign cfg_io_cfg_addr = io_cfg_addr[0]; // @[PE.scala 91:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 92:19]
endmodule
module GPE_28(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [3:0] alu_io_config; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 50:19]
  wire [31:0] alu_io_out; // @[PE.scala 50:19]
  wire  rf_clock; // @[PE.scala 51:18]
  wire  rf_reset; // @[PE.scala 51:18]
  wire  rf_io_en; // @[PE.scala 51:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 51:18]
  wire  DelayPipe_clock; // @[PE.scala 52:54]
  wire  DelayPipe_reset; // @[PE.scala 52:54]
  wire  DelayPipe_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 52:54]
  wire  DelayPipe_1_clock; // @[PE.scala 52:54]
  wire  DelayPipe_1_reset; // @[PE.scala 52:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 52:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 55:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 55:49]
  wire  cfg_clock; // @[PE.scala 89:19]
  wire  cfg_reset; // @[PE.scala 89:19]
  wire  cfg_io_cfg_en; // @[PE.scala 89:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 89:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 89:19]
  wire [47:0] cfg_io_out_0; // @[PE.scala 89:19]
  wire  _T_1 = 10'h56 == io_cfg_addr[11:2]; // @[PE.scala 90:48]
  wire [47:0] cfgOut = cfg_io_out_0; // @[PE.scala 96:20 PE.scala 97:10]
  ALU alu ( // @[PE.scala 50:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 51:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 52:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 52:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_16 Muxn ( // @[PE.scala 55:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_16 Muxn_1 ( // @[PE.scala 55:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_16 cfg ( // @[PE.scala 89:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 77:13]
  assign alu_io_config = cfgOut[35:32]; // @[PE.scala 100:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 71:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 71:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 75:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 76:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_io_config = cfgOut[38:36]; // @[PE.scala 113:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 70:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_1_io_config = cfgOut[41:39]; // @[PE.scala 113:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 70:23]
  assign Muxn_io_config = cfgOut[44:42]; // @[PE.scala 121:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 62:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 62:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 62:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 62:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign Muxn_1_io_config = cfgOut[47:45]; // @[PE.scala 121:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 62:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 62:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 62:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 62:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 90:17]
  assign cfg_io_cfg_addr = io_cfg_addr[0]; // @[PE.scala 91:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 92:19]
endmodule
module GPE_29(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [3:0] alu_io_config; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 50:19]
  wire [31:0] alu_io_out; // @[PE.scala 50:19]
  wire  rf_clock; // @[PE.scala 51:18]
  wire  rf_reset; // @[PE.scala 51:18]
  wire  rf_io_en; // @[PE.scala 51:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 51:18]
  wire  DelayPipe_clock; // @[PE.scala 52:54]
  wire  DelayPipe_reset; // @[PE.scala 52:54]
  wire  DelayPipe_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 52:54]
  wire  DelayPipe_1_clock; // @[PE.scala 52:54]
  wire  DelayPipe_1_reset; // @[PE.scala 52:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 52:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 55:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 55:49]
  wire  cfg_clock; // @[PE.scala 89:19]
  wire  cfg_reset; // @[PE.scala 89:19]
  wire  cfg_io_cfg_en; // @[PE.scala 89:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 89:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 89:19]
  wire [47:0] cfg_io_out_0; // @[PE.scala 89:19]
  wire  _T_1 = 10'h57 == io_cfg_addr[11:2]; // @[PE.scala 90:48]
  wire [47:0] cfgOut = cfg_io_out_0; // @[PE.scala 96:20 PE.scala 97:10]
  ALU alu ( // @[PE.scala 50:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 51:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 52:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 52:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_16 Muxn ( // @[PE.scala 55:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_16 Muxn_1 ( // @[PE.scala 55:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_16 cfg ( // @[PE.scala 89:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 77:13]
  assign alu_io_config = cfgOut[35:32]; // @[PE.scala 100:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 71:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 71:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 75:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 76:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_io_config = cfgOut[38:36]; // @[PE.scala 113:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 70:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_1_io_config = cfgOut[41:39]; // @[PE.scala 113:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 70:23]
  assign Muxn_io_config = cfgOut[44:42]; // @[PE.scala 121:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 62:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 62:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 62:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 62:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign Muxn_1_io_config = cfgOut[47:45]; // @[PE.scala 121:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 62:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 62:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 62:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 62:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 90:17]
  assign cfg_io_cfg_addr = io_cfg_addr[0]; // @[PE.scala 91:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 92:19]
endmodule
module GPE_30(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [3:0] alu_io_config; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 50:19]
  wire [31:0] alu_io_out; // @[PE.scala 50:19]
  wire  rf_clock; // @[PE.scala 51:18]
  wire  rf_reset; // @[PE.scala 51:18]
  wire  rf_io_en; // @[PE.scala 51:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 51:18]
  wire  DelayPipe_clock; // @[PE.scala 52:54]
  wire  DelayPipe_reset; // @[PE.scala 52:54]
  wire  DelayPipe_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 52:54]
  wire  DelayPipe_1_clock; // @[PE.scala 52:54]
  wire  DelayPipe_1_reset; // @[PE.scala 52:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 52:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 55:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 55:49]
  wire  cfg_clock; // @[PE.scala 89:19]
  wire  cfg_reset; // @[PE.scala 89:19]
  wire  cfg_io_cfg_en; // @[PE.scala 89:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 89:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 89:19]
  wire [47:0] cfg_io_out_0; // @[PE.scala 89:19]
  wire  _T_1 = 10'h58 == io_cfg_addr[11:2]; // @[PE.scala 90:48]
  wire [47:0] cfgOut = cfg_io_out_0; // @[PE.scala 96:20 PE.scala 97:10]
  ALU alu ( // @[PE.scala 50:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 51:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 52:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 52:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_16 Muxn ( // @[PE.scala 55:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_16 Muxn_1 ( // @[PE.scala 55:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_16 cfg ( // @[PE.scala 89:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 77:13]
  assign alu_io_config = cfgOut[35:32]; // @[PE.scala 100:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 71:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 71:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 75:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 76:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_io_config = cfgOut[38:36]; // @[PE.scala 113:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 70:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_1_io_config = cfgOut[41:39]; // @[PE.scala 113:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 70:23]
  assign Muxn_io_config = cfgOut[44:42]; // @[PE.scala 121:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 62:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 62:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 62:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 62:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign Muxn_1_io_config = cfgOut[47:45]; // @[PE.scala 121:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 62:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 62:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 62:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 62:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 90:17]
  assign cfg_io_cfg_addr = io_cfg_addr[0]; // @[PE.scala 91:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 92:19]
endmodule
module GPE_31(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [3:0] alu_io_config; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 50:19]
  wire [31:0] alu_io_out; // @[PE.scala 50:19]
  wire  rf_clock; // @[PE.scala 51:18]
  wire  rf_reset; // @[PE.scala 51:18]
  wire  rf_io_en; // @[PE.scala 51:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 51:18]
  wire  DelayPipe_clock; // @[PE.scala 52:54]
  wire  DelayPipe_reset; // @[PE.scala 52:54]
  wire  DelayPipe_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 52:54]
  wire  DelayPipe_1_clock; // @[PE.scala 52:54]
  wire  DelayPipe_1_reset; // @[PE.scala 52:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 52:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 55:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 55:49]
  wire  cfg_clock; // @[PE.scala 89:19]
  wire  cfg_reset; // @[PE.scala 89:19]
  wire  cfg_io_cfg_en; // @[PE.scala 89:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 89:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 89:19]
  wire [47:0] cfg_io_out_0; // @[PE.scala 89:19]
  wire  _T_1 = 10'h59 == io_cfg_addr[11:2]; // @[PE.scala 90:48]
  wire [47:0] cfgOut = cfg_io_out_0; // @[PE.scala 96:20 PE.scala 97:10]
  ALU alu ( // @[PE.scala 50:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 51:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 52:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 52:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_16 Muxn ( // @[PE.scala 55:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_16 Muxn_1 ( // @[PE.scala 55:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_16 cfg ( // @[PE.scala 89:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 77:13]
  assign alu_io_config = cfgOut[35:32]; // @[PE.scala 100:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 71:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 71:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 75:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 76:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_io_config = cfgOut[38:36]; // @[PE.scala 113:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 70:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_1_io_config = cfgOut[41:39]; // @[PE.scala 113:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 70:23]
  assign Muxn_io_config = cfgOut[44:42]; // @[PE.scala 121:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 62:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 62:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 62:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 62:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign Muxn_1_io_config = cfgOut[47:45]; // @[PE.scala 121:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 62:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 62:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 62:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 62:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 90:17]
  assign cfg_io_cfg_addr = io_cfg_addr[0]; // @[PE.scala 91:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 92:19]
endmodule
module GPE_32(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [3:0] alu_io_config; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 50:19]
  wire [31:0] alu_io_out; // @[PE.scala 50:19]
  wire  rf_clock; // @[PE.scala 51:18]
  wire  rf_reset; // @[PE.scala 51:18]
  wire  rf_io_en; // @[PE.scala 51:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 51:18]
  wire  DelayPipe_clock; // @[PE.scala 52:54]
  wire  DelayPipe_reset; // @[PE.scala 52:54]
  wire  DelayPipe_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 52:54]
  wire  DelayPipe_1_clock; // @[PE.scala 52:54]
  wire  DelayPipe_1_reset; // @[PE.scala 52:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 52:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 55:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 55:49]
  wire  cfg_clock; // @[PE.scala 89:19]
  wire  cfg_reset; // @[PE.scala 89:19]
  wire  cfg_io_cfg_en; // @[PE.scala 89:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 89:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 89:19]
  wire [47:0] cfg_io_out_0; // @[PE.scala 89:19]
  wire  _T_1 = 10'h64 == io_cfg_addr[11:2]; // @[PE.scala 90:48]
  wire [47:0] cfgOut = cfg_io_out_0; // @[PE.scala 96:20 PE.scala 97:10]
  ALU alu ( // @[PE.scala 50:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 51:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 52:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 52:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_16 Muxn ( // @[PE.scala 55:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_16 Muxn_1 ( // @[PE.scala 55:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_16 cfg ( // @[PE.scala 89:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 77:13]
  assign alu_io_config = cfgOut[35:32]; // @[PE.scala 100:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 71:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 71:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 75:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 76:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_io_config = cfgOut[38:36]; // @[PE.scala 113:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 70:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_1_io_config = cfgOut[41:39]; // @[PE.scala 113:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 70:23]
  assign Muxn_io_config = cfgOut[44:42]; // @[PE.scala 121:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 62:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 62:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 62:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 62:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign Muxn_1_io_config = cfgOut[47:45]; // @[PE.scala 121:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 62:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 62:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 62:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 62:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 90:17]
  assign cfg_io_cfg_addr = io_cfg_addr[0]; // @[PE.scala 91:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 92:19]
endmodule
module GPE_33(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [3:0] alu_io_config; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 50:19]
  wire [31:0] alu_io_out; // @[PE.scala 50:19]
  wire  rf_clock; // @[PE.scala 51:18]
  wire  rf_reset; // @[PE.scala 51:18]
  wire  rf_io_en; // @[PE.scala 51:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 51:18]
  wire  DelayPipe_clock; // @[PE.scala 52:54]
  wire  DelayPipe_reset; // @[PE.scala 52:54]
  wire  DelayPipe_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 52:54]
  wire  DelayPipe_1_clock; // @[PE.scala 52:54]
  wire  DelayPipe_1_reset; // @[PE.scala 52:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 52:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 55:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 55:49]
  wire  cfg_clock; // @[PE.scala 89:19]
  wire  cfg_reset; // @[PE.scala 89:19]
  wire  cfg_io_cfg_en; // @[PE.scala 89:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 89:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 89:19]
  wire [47:0] cfg_io_out_0; // @[PE.scala 89:19]
  wire  _T_1 = 10'h65 == io_cfg_addr[11:2]; // @[PE.scala 90:48]
  wire [47:0] cfgOut = cfg_io_out_0; // @[PE.scala 96:20 PE.scala 97:10]
  ALU alu ( // @[PE.scala 50:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 51:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 52:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 52:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_16 Muxn ( // @[PE.scala 55:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_16 Muxn_1 ( // @[PE.scala 55:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_16 cfg ( // @[PE.scala 89:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 77:13]
  assign alu_io_config = cfgOut[35:32]; // @[PE.scala 100:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 71:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 71:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 75:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 76:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_io_config = cfgOut[38:36]; // @[PE.scala 113:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 70:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_1_io_config = cfgOut[41:39]; // @[PE.scala 113:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 70:23]
  assign Muxn_io_config = cfgOut[44:42]; // @[PE.scala 121:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 62:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 62:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 62:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 62:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign Muxn_1_io_config = cfgOut[47:45]; // @[PE.scala 121:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 62:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 62:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 62:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 62:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 90:17]
  assign cfg_io_cfg_addr = io_cfg_addr[0]; // @[PE.scala 91:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 92:19]
endmodule
module GPE_34(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [3:0] alu_io_config; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 50:19]
  wire [31:0] alu_io_out; // @[PE.scala 50:19]
  wire  rf_clock; // @[PE.scala 51:18]
  wire  rf_reset; // @[PE.scala 51:18]
  wire  rf_io_en; // @[PE.scala 51:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 51:18]
  wire  DelayPipe_clock; // @[PE.scala 52:54]
  wire  DelayPipe_reset; // @[PE.scala 52:54]
  wire  DelayPipe_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 52:54]
  wire  DelayPipe_1_clock; // @[PE.scala 52:54]
  wire  DelayPipe_1_reset; // @[PE.scala 52:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 52:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 55:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 55:49]
  wire  cfg_clock; // @[PE.scala 89:19]
  wire  cfg_reset; // @[PE.scala 89:19]
  wire  cfg_io_cfg_en; // @[PE.scala 89:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 89:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 89:19]
  wire [47:0] cfg_io_out_0; // @[PE.scala 89:19]
  wire  _T_1 = 10'h66 == io_cfg_addr[11:2]; // @[PE.scala 90:48]
  wire [47:0] cfgOut = cfg_io_out_0; // @[PE.scala 96:20 PE.scala 97:10]
  ALU alu ( // @[PE.scala 50:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 51:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 52:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 52:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_16 Muxn ( // @[PE.scala 55:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_16 Muxn_1 ( // @[PE.scala 55:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_16 cfg ( // @[PE.scala 89:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 77:13]
  assign alu_io_config = cfgOut[35:32]; // @[PE.scala 100:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 71:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 71:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 75:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 76:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_io_config = cfgOut[38:36]; // @[PE.scala 113:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 70:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_1_io_config = cfgOut[41:39]; // @[PE.scala 113:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 70:23]
  assign Muxn_io_config = cfgOut[44:42]; // @[PE.scala 121:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 62:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 62:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 62:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 62:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign Muxn_1_io_config = cfgOut[47:45]; // @[PE.scala 121:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 62:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 62:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 62:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 62:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 90:17]
  assign cfg_io_cfg_addr = io_cfg_addr[0]; // @[PE.scala 91:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 92:19]
endmodule
module GPE_35(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [3:0] alu_io_config; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 50:19]
  wire [31:0] alu_io_out; // @[PE.scala 50:19]
  wire  rf_clock; // @[PE.scala 51:18]
  wire  rf_reset; // @[PE.scala 51:18]
  wire  rf_io_en; // @[PE.scala 51:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 51:18]
  wire  DelayPipe_clock; // @[PE.scala 52:54]
  wire  DelayPipe_reset; // @[PE.scala 52:54]
  wire  DelayPipe_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 52:54]
  wire  DelayPipe_1_clock; // @[PE.scala 52:54]
  wire  DelayPipe_1_reset; // @[PE.scala 52:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 52:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 55:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 55:49]
  wire  cfg_clock; // @[PE.scala 89:19]
  wire  cfg_reset; // @[PE.scala 89:19]
  wire  cfg_io_cfg_en; // @[PE.scala 89:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 89:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 89:19]
  wire [47:0] cfg_io_out_0; // @[PE.scala 89:19]
  wire  _T_1 = 10'h67 == io_cfg_addr[11:2]; // @[PE.scala 90:48]
  wire [47:0] cfgOut = cfg_io_out_0; // @[PE.scala 96:20 PE.scala 97:10]
  ALU alu ( // @[PE.scala 50:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 51:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 52:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 52:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_16 Muxn ( // @[PE.scala 55:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_16 Muxn_1 ( // @[PE.scala 55:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_16 cfg ( // @[PE.scala 89:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 77:13]
  assign alu_io_config = cfgOut[35:32]; // @[PE.scala 100:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 71:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 71:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 75:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 76:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_io_config = cfgOut[38:36]; // @[PE.scala 113:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 70:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_1_io_config = cfgOut[41:39]; // @[PE.scala 113:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 70:23]
  assign Muxn_io_config = cfgOut[44:42]; // @[PE.scala 121:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 62:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 62:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 62:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 62:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign Muxn_1_io_config = cfgOut[47:45]; // @[PE.scala 121:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 62:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 62:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 62:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 62:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 90:17]
  assign cfg_io_cfg_addr = io_cfg_addr[0]; // @[PE.scala 91:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 92:19]
endmodule
module GPE_36(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [3:0] alu_io_config; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 50:19]
  wire [31:0] alu_io_out; // @[PE.scala 50:19]
  wire  rf_clock; // @[PE.scala 51:18]
  wire  rf_reset; // @[PE.scala 51:18]
  wire  rf_io_en; // @[PE.scala 51:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 51:18]
  wire  DelayPipe_clock; // @[PE.scala 52:54]
  wire  DelayPipe_reset; // @[PE.scala 52:54]
  wire  DelayPipe_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 52:54]
  wire  DelayPipe_1_clock; // @[PE.scala 52:54]
  wire  DelayPipe_1_reset; // @[PE.scala 52:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 52:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 55:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 55:49]
  wire  cfg_clock; // @[PE.scala 89:19]
  wire  cfg_reset; // @[PE.scala 89:19]
  wire  cfg_io_cfg_en; // @[PE.scala 89:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 89:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 89:19]
  wire [47:0] cfg_io_out_0; // @[PE.scala 89:19]
  wire  _T_1 = 10'h68 == io_cfg_addr[11:2]; // @[PE.scala 90:48]
  wire [47:0] cfgOut = cfg_io_out_0; // @[PE.scala 96:20 PE.scala 97:10]
  ALU alu ( // @[PE.scala 50:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 51:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 52:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 52:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_16 Muxn ( // @[PE.scala 55:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_16 Muxn_1 ( // @[PE.scala 55:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_16 cfg ( // @[PE.scala 89:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 77:13]
  assign alu_io_config = cfgOut[35:32]; // @[PE.scala 100:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 71:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 71:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 75:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 76:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_io_config = cfgOut[38:36]; // @[PE.scala 113:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 70:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_1_io_config = cfgOut[41:39]; // @[PE.scala 113:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 70:23]
  assign Muxn_io_config = cfgOut[44:42]; // @[PE.scala 121:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 62:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 62:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 62:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 62:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign Muxn_1_io_config = cfgOut[47:45]; // @[PE.scala 121:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 62:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 62:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 62:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 62:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 90:17]
  assign cfg_io_cfg_addr = io_cfg_addr[0]; // @[PE.scala 91:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 92:19]
endmodule
module GPE_37(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [3:0] alu_io_config; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 50:19]
  wire [31:0] alu_io_out; // @[PE.scala 50:19]
  wire  rf_clock; // @[PE.scala 51:18]
  wire  rf_reset; // @[PE.scala 51:18]
  wire  rf_io_en; // @[PE.scala 51:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 51:18]
  wire  DelayPipe_clock; // @[PE.scala 52:54]
  wire  DelayPipe_reset; // @[PE.scala 52:54]
  wire  DelayPipe_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 52:54]
  wire  DelayPipe_1_clock; // @[PE.scala 52:54]
  wire  DelayPipe_1_reset; // @[PE.scala 52:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 52:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 55:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 55:49]
  wire  cfg_clock; // @[PE.scala 89:19]
  wire  cfg_reset; // @[PE.scala 89:19]
  wire  cfg_io_cfg_en; // @[PE.scala 89:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 89:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 89:19]
  wire [47:0] cfg_io_out_0; // @[PE.scala 89:19]
  wire  _T_1 = 10'h69 == io_cfg_addr[11:2]; // @[PE.scala 90:48]
  wire [47:0] cfgOut = cfg_io_out_0; // @[PE.scala 96:20 PE.scala 97:10]
  ALU alu ( // @[PE.scala 50:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 51:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 52:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 52:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_16 Muxn ( // @[PE.scala 55:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_16 Muxn_1 ( // @[PE.scala 55:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_16 cfg ( // @[PE.scala 89:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 77:13]
  assign alu_io_config = cfgOut[35:32]; // @[PE.scala 100:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 71:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 71:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 75:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 76:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_io_config = cfgOut[38:36]; // @[PE.scala 113:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 70:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_1_io_config = cfgOut[41:39]; // @[PE.scala 113:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 70:23]
  assign Muxn_io_config = cfgOut[44:42]; // @[PE.scala 121:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 62:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 62:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 62:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 62:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign Muxn_1_io_config = cfgOut[47:45]; // @[PE.scala 121:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 62:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 62:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 62:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 62:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 90:17]
  assign cfg_io_cfg_addr = io_cfg_addr[0]; // @[PE.scala 91:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 92:19]
endmodule
module GPE_38(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [3:0] alu_io_config; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 50:19]
  wire [31:0] alu_io_out; // @[PE.scala 50:19]
  wire  rf_clock; // @[PE.scala 51:18]
  wire  rf_reset; // @[PE.scala 51:18]
  wire  rf_io_en; // @[PE.scala 51:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 51:18]
  wire  DelayPipe_clock; // @[PE.scala 52:54]
  wire  DelayPipe_reset; // @[PE.scala 52:54]
  wire  DelayPipe_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 52:54]
  wire  DelayPipe_1_clock; // @[PE.scala 52:54]
  wire  DelayPipe_1_reset; // @[PE.scala 52:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 52:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 55:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 55:49]
  wire  cfg_clock; // @[PE.scala 89:19]
  wire  cfg_reset; // @[PE.scala 89:19]
  wire  cfg_io_cfg_en; // @[PE.scala 89:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 89:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 89:19]
  wire [47:0] cfg_io_out_0; // @[PE.scala 89:19]
  wire  _T_1 = 10'h6a == io_cfg_addr[11:2]; // @[PE.scala 90:48]
  wire [47:0] cfgOut = cfg_io_out_0; // @[PE.scala 96:20 PE.scala 97:10]
  ALU alu ( // @[PE.scala 50:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 51:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 52:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 52:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_16 Muxn ( // @[PE.scala 55:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_16 Muxn_1 ( // @[PE.scala 55:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_16 cfg ( // @[PE.scala 89:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 77:13]
  assign alu_io_config = cfgOut[35:32]; // @[PE.scala 100:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 71:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 71:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 75:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 76:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_io_config = cfgOut[38:36]; // @[PE.scala 113:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 70:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_1_io_config = cfgOut[41:39]; // @[PE.scala 113:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 70:23]
  assign Muxn_io_config = cfgOut[44:42]; // @[PE.scala 121:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 62:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 62:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 62:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 62:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign Muxn_1_io_config = cfgOut[47:45]; // @[PE.scala 121:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 62:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 62:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 62:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 62:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 90:17]
  assign cfg_io_cfg_addr = io_cfg_addr[0]; // @[PE.scala 91:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 92:19]
endmodule
module GPE_39(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [3:0] alu_io_config; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 50:19]
  wire [31:0] alu_io_out; // @[PE.scala 50:19]
  wire  rf_clock; // @[PE.scala 51:18]
  wire  rf_reset; // @[PE.scala 51:18]
  wire  rf_io_en; // @[PE.scala 51:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 51:18]
  wire  DelayPipe_clock; // @[PE.scala 52:54]
  wire  DelayPipe_reset; // @[PE.scala 52:54]
  wire  DelayPipe_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 52:54]
  wire  DelayPipe_1_clock; // @[PE.scala 52:54]
  wire  DelayPipe_1_reset; // @[PE.scala 52:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 52:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 55:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 55:49]
  wire  cfg_clock; // @[PE.scala 89:19]
  wire  cfg_reset; // @[PE.scala 89:19]
  wire  cfg_io_cfg_en; // @[PE.scala 89:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 89:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 89:19]
  wire [47:0] cfg_io_out_0; // @[PE.scala 89:19]
  wire  _T_1 = 10'h6b == io_cfg_addr[11:2]; // @[PE.scala 90:48]
  wire [47:0] cfgOut = cfg_io_out_0; // @[PE.scala 96:20 PE.scala 97:10]
  ALU alu ( // @[PE.scala 50:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 51:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 52:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 52:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_16 Muxn ( // @[PE.scala 55:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_16 Muxn_1 ( // @[PE.scala 55:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_16 cfg ( // @[PE.scala 89:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 77:13]
  assign alu_io_config = cfgOut[35:32]; // @[PE.scala 100:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 71:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 71:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 75:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 76:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_io_config = cfgOut[38:36]; // @[PE.scala 113:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 70:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_1_io_config = cfgOut[41:39]; // @[PE.scala 113:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 70:23]
  assign Muxn_io_config = cfgOut[44:42]; // @[PE.scala 121:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 62:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 62:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 62:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 62:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign Muxn_1_io_config = cfgOut[47:45]; // @[PE.scala 121:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 62:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 62:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 62:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 62:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 90:17]
  assign cfg_io_cfg_addr = io_cfg_addr[0]; // @[PE.scala 91:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 92:19]
endmodule
module GPE_40(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [3:0] alu_io_config; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 50:19]
  wire [31:0] alu_io_out; // @[PE.scala 50:19]
  wire  rf_clock; // @[PE.scala 51:18]
  wire  rf_reset; // @[PE.scala 51:18]
  wire  rf_io_en; // @[PE.scala 51:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 51:18]
  wire  DelayPipe_clock; // @[PE.scala 52:54]
  wire  DelayPipe_reset; // @[PE.scala 52:54]
  wire  DelayPipe_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 52:54]
  wire  DelayPipe_1_clock; // @[PE.scala 52:54]
  wire  DelayPipe_1_reset; // @[PE.scala 52:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 52:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 55:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 55:49]
  wire  cfg_clock; // @[PE.scala 89:19]
  wire  cfg_reset; // @[PE.scala 89:19]
  wire  cfg_io_cfg_en; // @[PE.scala 89:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 89:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 89:19]
  wire [47:0] cfg_io_out_0; // @[PE.scala 89:19]
  wire  _T_1 = 10'h76 == io_cfg_addr[11:2]; // @[PE.scala 90:48]
  wire [47:0] cfgOut = cfg_io_out_0; // @[PE.scala 96:20 PE.scala 97:10]
  ALU alu ( // @[PE.scala 50:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 51:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 52:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 52:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_16 Muxn ( // @[PE.scala 55:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_16 Muxn_1 ( // @[PE.scala 55:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_16 cfg ( // @[PE.scala 89:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 77:13]
  assign alu_io_config = cfgOut[35:32]; // @[PE.scala 100:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 71:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 71:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 75:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 76:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_io_config = cfgOut[38:36]; // @[PE.scala 113:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 70:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_1_io_config = cfgOut[41:39]; // @[PE.scala 113:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 70:23]
  assign Muxn_io_config = cfgOut[44:42]; // @[PE.scala 121:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 62:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 62:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 62:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 62:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign Muxn_1_io_config = cfgOut[47:45]; // @[PE.scala 121:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 62:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 62:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 62:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 62:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 90:17]
  assign cfg_io_cfg_addr = io_cfg_addr[0]; // @[PE.scala 91:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 92:19]
endmodule
module GPE_41(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [3:0] alu_io_config; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 50:19]
  wire [31:0] alu_io_out; // @[PE.scala 50:19]
  wire  rf_clock; // @[PE.scala 51:18]
  wire  rf_reset; // @[PE.scala 51:18]
  wire  rf_io_en; // @[PE.scala 51:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 51:18]
  wire  DelayPipe_clock; // @[PE.scala 52:54]
  wire  DelayPipe_reset; // @[PE.scala 52:54]
  wire  DelayPipe_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 52:54]
  wire  DelayPipe_1_clock; // @[PE.scala 52:54]
  wire  DelayPipe_1_reset; // @[PE.scala 52:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 52:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 55:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 55:49]
  wire  cfg_clock; // @[PE.scala 89:19]
  wire  cfg_reset; // @[PE.scala 89:19]
  wire  cfg_io_cfg_en; // @[PE.scala 89:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 89:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 89:19]
  wire [47:0] cfg_io_out_0; // @[PE.scala 89:19]
  wire  _T_1 = 10'h77 == io_cfg_addr[11:2]; // @[PE.scala 90:48]
  wire [47:0] cfgOut = cfg_io_out_0; // @[PE.scala 96:20 PE.scala 97:10]
  ALU alu ( // @[PE.scala 50:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 51:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 52:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 52:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_16 Muxn ( // @[PE.scala 55:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_16 Muxn_1 ( // @[PE.scala 55:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_16 cfg ( // @[PE.scala 89:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 77:13]
  assign alu_io_config = cfgOut[35:32]; // @[PE.scala 100:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 71:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 71:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 75:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 76:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_io_config = cfgOut[38:36]; // @[PE.scala 113:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 70:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_1_io_config = cfgOut[41:39]; // @[PE.scala 113:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 70:23]
  assign Muxn_io_config = cfgOut[44:42]; // @[PE.scala 121:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 62:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 62:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 62:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 62:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign Muxn_1_io_config = cfgOut[47:45]; // @[PE.scala 121:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 62:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 62:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 62:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 62:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 90:17]
  assign cfg_io_cfg_addr = io_cfg_addr[0]; // @[PE.scala 91:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 92:19]
endmodule
module GPE_42(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [3:0] alu_io_config; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 50:19]
  wire [31:0] alu_io_out; // @[PE.scala 50:19]
  wire  rf_clock; // @[PE.scala 51:18]
  wire  rf_reset; // @[PE.scala 51:18]
  wire  rf_io_en; // @[PE.scala 51:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 51:18]
  wire  DelayPipe_clock; // @[PE.scala 52:54]
  wire  DelayPipe_reset; // @[PE.scala 52:54]
  wire  DelayPipe_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 52:54]
  wire  DelayPipe_1_clock; // @[PE.scala 52:54]
  wire  DelayPipe_1_reset; // @[PE.scala 52:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 52:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 55:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 55:49]
  wire  cfg_clock; // @[PE.scala 89:19]
  wire  cfg_reset; // @[PE.scala 89:19]
  wire  cfg_io_cfg_en; // @[PE.scala 89:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 89:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 89:19]
  wire [47:0] cfg_io_out_0; // @[PE.scala 89:19]
  wire  _T_1 = 10'h78 == io_cfg_addr[11:2]; // @[PE.scala 90:48]
  wire [47:0] cfgOut = cfg_io_out_0; // @[PE.scala 96:20 PE.scala 97:10]
  ALU alu ( // @[PE.scala 50:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 51:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 52:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 52:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_16 Muxn ( // @[PE.scala 55:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_16 Muxn_1 ( // @[PE.scala 55:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_16 cfg ( // @[PE.scala 89:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 77:13]
  assign alu_io_config = cfgOut[35:32]; // @[PE.scala 100:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 71:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 71:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 75:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 76:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_io_config = cfgOut[38:36]; // @[PE.scala 113:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 70:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_1_io_config = cfgOut[41:39]; // @[PE.scala 113:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 70:23]
  assign Muxn_io_config = cfgOut[44:42]; // @[PE.scala 121:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 62:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 62:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 62:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 62:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign Muxn_1_io_config = cfgOut[47:45]; // @[PE.scala 121:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 62:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 62:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 62:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 62:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 90:17]
  assign cfg_io_cfg_addr = io_cfg_addr[0]; // @[PE.scala 91:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 92:19]
endmodule
module GPE_43(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [3:0] alu_io_config; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 50:19]
  wire [31:0] alu_io_out; // @[PE.scala 50:19]
  wire  rf_clock; // @[PE.scala 51:18]
  wire  rf_reset; // @[PE.scala 51:18]
  wire  rf_io_en; // @[PE.scala 51:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 51:18]
  wire  DelayPipe_clock; // @[PE.scala 52:54]
  wire  DelayPipe_reset; // @[PE.scala 52:54]
  wire  DelayPipe_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 52:54]
  wire  DelayPipe_1_clock; // @[PE.scala 52:54]
  wire  DelayPipe_1_reset; // @[PE.scala 52:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 52:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 55:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 55:49]
  wire  cfg_clock; // @[PE.scala 89:19]
  wire  cfg_reset; // @[PE.scala 89:19]
  wire  cfg_io_cfg_en; // @[PE.scala 89:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 89:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 89:19]
  wire [47:0] cfg_io_out_0; // @[PE.scala 89:19]
  wire  _T_1 = 10'h79 == io_cfg_addr[11:2]; // @[PE.scala 90:48]
  wire [47:0] cfgOut = cfg_io_out_0; // @[PE.scala 96:20 PE.scala 97:10]
  ALU alu ( // @[PE.scala 50:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 51:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 52:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 52:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_16 Muxn ( // @[PE.scala 55:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_16 Muxn_1 ( // @[PE.scala 55:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_16 cfg ( // @[PE.scala 89:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 77:13]
  assign alu_io_config = cfgOut[35:32]; // @[PE.scala 100:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 71:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 71:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 75:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 76:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_io_config = cfgOut[38:36]; // @[PE.scala 113:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 70:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_1_io_config = cfgOut[41:39]; // @[PE.scala 113:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 70:23]
  assign Muxn_io_config = cfgOut[44:42]; // @[PE.scala 121:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 62:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 62:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 62:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 62:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign Muxn_1_io_config = cfgOut[47:45]; // @[PE.scala 121:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 62:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 62:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 62:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 62:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 90:17]
  assign cfg_io_cfg_addr = io_cfg_addr[0]; // @[PE.scala 91:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 92:19]
endmodule
module GPE_44(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [3:0] alu_io_config; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 50:19]
  wire [31:0] alu_io_out; // @[PE.scala 50:19]
  wire  rf_clock; // @[PE.scala 51:18]
  wire  rf_reset; // @[PE.scala 51:18]
  wire  rf_io_en; // @[PE.scala 51:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 51:18]
  wire  DelayPipe_clock; // @[PE.scala 52:54]
  wire  DelayPipe_reset; // @[PE.scala 52:54]
  wire  DelayPipe_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 52:54]
  wire  DelayPipe_1_clock; // @[PE.scala 52:54]
  wire  DelayPipe_1_reset; // @[PE.scala 52:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 52:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 55:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 55:49]
  wire  cfg_clock; // @[PE.scala 89:19]
  wire  cfg_reset; // @[PE.scala 89:19]
  wire  cfg_io_cfg_en; // @[PE.scala 89:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 89:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 89:19]
  wire [47:0] cfg_io_out_0; // @[PE.scala 89:19]
  wire  _T_1 = 10'h7a == io_cfg_addr[11:2]; // @[PE.scala 90:48]
  wire [47:0] cfgOut = cfg_io_out_0; // @[PE.scala 96:20 PE.scala 97:10]
  ALU alu ( // @[PE.scala 50:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 51:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 52:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 52:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_16 Muxn ( // @[PE.scala 55:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_16 Muxn_1 ( // @[PE.scala 55:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_16 cfg ( // @[PE.scala 89:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 77:13]
  assign alu_io_config = cfgOut[35:32]; // @[PE.scala 100:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 71:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 71:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 75:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 76:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_io_config = cfgOut[38:36]; // @[PE.scala 113:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 70:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_1_io_config = cfgOut[41:39]; // @[PE.scala 113:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 70:23]
  assign Muxn_io_config = cfgOut[44:42]; // @[PE.scala 121:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 62:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 62:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 62:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 62:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign Muxn_1_io_config = cfgOut[47:45]; // @[PE.scala 121:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 62:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 62:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 62:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 62:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 90:17]
  assign cfg_io_cfg_addr = io_cfg_addr[0]; // @[PE.scala 91:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 92:19]
endmodule
module GPE_45(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [3:0] alu_io_config; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 50:19]
  wire [31:0] alu_io_out; // @[PE.scala 50:19]
  wire  rf_clock; // @[PE.scala 51:18]
  wire  rf_reset; // @[PE.scala 51:18]
  wire  rf_io_en; // @[PE.scala 51:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 51:18]
  wire  DelayPipe_clock; // @[PE.scala 52:54]
  wire  DelayPipe_reset; // @[PE.scala 52:54]
  wire  DelayPipe_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 52:54]
  wire  DelayPipe_1_clock; // @[PE.scala 52:54]
  wire  DelayPipe_1_reset; // @[PE.scala 52:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 52:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 55:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 55:49]
  wire  cfg_clock; // @[PE.scala 89:19]
  wire  cfg_reset; // @[PE.scala 89:19]
  wire  cfg_io_cfg_en; // @[PE.scala 89:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 89:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 89:19]
  wire [47:0] cfg_io_out_0; // @[PE.scala 89:19]
  wire  _T_1 = 10'h7b == io_cfg_addr[11:2]; // @[PE.scala 90:48]
  wire [47:0] cfgOut = cfg_io_out_0; // @[PE.scala 96:20 PE.scala 97:10]
  ALU alu ( // @[PE.scala 50:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 51:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 52:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 52:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_16 Muxn ( // @[PE.scala 55:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_16 Muxn_1 ( // @[PE.scala 55:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_16 cfg ( // @[PE.scala 89:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 77:13]
  assign alu_io_config = cfgOut[35:32]; // @[PE.scala 100:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 71:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 71:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 75:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 76:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_io_config = cfgOut[38:36]; // @[PE.scala 113:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 70:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_1_io_config = cfgOut[41:39]; // @[PE.scala 113:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 70:23]
  assign Muxn_io_config = cfgOut[44:42]; // @[PE.scala 121:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 62:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 62:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 62:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 62:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign Muxn_1_io_config = cfgOut[47:45]; // @[PE.scala 121:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 62:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 62:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 62:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 62:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 90:17]
  assign cfg_io_cfg_addr = io_cfg_addr[0]; // @[PE.scala 91:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 92:19]
endmodule
module GPE_46(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [3:0] alu_io_config; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 50:19]
  wire [31:0] alu_io_out; // @[PE.scala 50:19]
  wire  rf_clock; // @[PE.scala 51:18]
  wire  rf_reset; // @[PE.scala 51:18]
  wire  rf_io_en; // @[PE.scala 51:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 51:18]
  wire  DelayPipe_clock; // @[PE.scala 52:54]
  wire  DelayPipe_reset; // @[PE.scala 52:54]
  wire  DelayPipe_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 52:54]
  wire  DelayPipe_1_clock; // @[PE.scala 52:54]
  wire  DelayPipe_1_reset; // @[PE.scala 52:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 52:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 55:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 55:49]
  wire  cfg_clock; // @[PE.scala 89:19]
  wire  cfg_reset; // @[PE.scala 89:19]
  wire  cfg_io_cfg_en; // @[PE.scala 89:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 89:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 89:19]
  wire [47:0] cfg_io_out_0; // @[PE.scala 89:19]
  wire  _T_1 = 10'h7c == io_cfg_addr[11:2]; // @[PE.scala 90:48]
  wire [47:0] cfgOut = cfg_io_out_0; // @[PE.scala 96:20 PE.scala 97:10]
  ALU alu ( // @[PE.scala 50:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 51:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 52:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 52:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_16 Muxn ( // @[PE.scala 55:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_16 Muxn_1 ( // @[PE.scala 55:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_16 cfg ( // @[PE.scala 89:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 77:13]
  assign alu_io_config = cfgOut[35:32]; // @[PE.scala 100:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 71:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 71:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 75:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 76:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_io_config = cfgOut[38:36]; // @[PE.scala 113:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 70:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_1_io_config = cfgOut[41:39]; // @[PE.scala 113:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 70:23]
  assign Muxn_io_config = cfgOut[44:42]; // @[PE.scala 121:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 62:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 62:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 62:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 62:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign Muxn_1_io_config = cfgOut[47:45]; // @[PE.scala 121:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 62:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 62:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 62:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 62:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 90:17]
  assign cfg_io_cfg_addr = io_cfg_addr[0]; // @[PE.scala 91:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 92:19]
endmodule
module GPE_47(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [3:0] alu_io_config; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 50:19]
  wire [31:0] alu_io_out; // @[PE.scala 50:19]
  wire  rf_clock; // @[PE.scala 51:18]
  wire  rf_reset; // @[PE.scala 51:18]
  wire  rf_io_en; // @[PE.scala 51:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 51:18]
  wire  DelayPipe_clock; // @[PE.scala 52:54]
  wire  DelayPipe_reset; // @[PE.scala 52:54]
  wire  DelayPipe_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 52:54]
  wire  DelayPipe_1_clock; // @[PE.scala 52:54]
  wire  DelayPipe_1_reset; // @[PE.scala 52:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 52:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 55:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 55:49]
  wire  cfg_clock; // @[PE.scala 89:19]
  wire  cfg_reset; // @[PE.scala 89:19]
  wire  cfg_io_cfg_en; // @[PE.scala 89:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 89:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 89:19]
  wire [47:0] cfg_io_out_0; // @[PE.scala 89:19]
  wire  _T_1 = 10'h7d == io_cfg_addr[11:2]; // @[PE.scala 90:48]
  wire [47:0] cfgOut = cfg_io_out_0; // @[PE.scala 96:20 PE.scala 97:10]
  ALU alu ( // @[PE.scala 50:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 51:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 52:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 52:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_16 Muxn ( // @[PE.scala 55:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_16 Muxn_1 ( // @[PE.scala 55:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_16 cfg ( // @[PE.scala 89:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 77:13]
  assign alu_io_config = cfgOut[35:32]; // @[PE.scala 100:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 71:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 71:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 75:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 76:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_io_config = cfgOut[38:36]; // @[PE.scala 113:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 70:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_1_io_config = cfgOut[41:39]; // @[PE.scala 113:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 70:23]
  assign Muxn_io_config = cfgOut[44:42]; // @[PE.scala 121:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 62:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 62:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 62:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 62:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign Muxn_1_io_config = cfgOut[47:45]; // @[PE.scala 121:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 62:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 62:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 62:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 62:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 90:17]
  assign cfg_io_cfg_addr = io_cfg_addr[0]; // @[PE.scala 91:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 92:19]
endmodule
module GPE_48(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [3:0] alu_io_config; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 50:19]
  wire [31:0] alu_io_out; // @[PE.scala 50:19]
  wire  rf_clock; // @[PE.scala 51:18]
  wire  rf_reset; // @[PE.scala 51:18]
  wire  rf_io_en; // @[PE.scala 51:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 51:18]
  wire  DelayPipe_clock; // @[PE.scala 52:54]
  wire  DelayPipe_reset; // @[PE.scala 52:54]
  wire  DelayPipe_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 52:54]
  wire  DelayPipe_1_clock; // @[PE.scala 52:54]
  wire  DelayPipe_1_reset; // @[PE.scala 52:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 52:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 55:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 55:49]
  wire  cfg_clock; // @[PE.scala 89:19]
  wire  cfg_reset; // @[PE.scala 89:19]
  wire  cfg_io_cfg_en; // @[PE.scala 89:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 89:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 89:19]
  wire [47:0] cfg_io_out_0; // @[PE.scala 89:19]
  wire  _T_1 = 10'h88 == io_cfg_addr[11:2]; // @[PE.scala 90:48]
  wire [47:0] cfgOut = cfg_io_out_0; // @[PE.scala 96:20 PE.scala 97:10]
  ALU alu ( // @[PE.scala 50:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 51:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 52:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 52:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_16 Muxn ( // @[PE.scala 55:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_16 Muxn_1 ( // @[PE.scala 55:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_16 cfg ( // @[PE.scala 89:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 77:13]
  assign alu_io_config = cfgOut[35:32]; // @[PE.scala 100:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 71:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 71:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 75:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 76:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_io_config = cfgOut[38:36]; // @[PE.scala 113:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 70:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_1_io_config = cfgOut[41:39]; // @[PE.scala 113:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 70:23]
  assign Muxn_io_config = cfgOut[44:42]; // @[PE.scala 121:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 62:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 62:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 62:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 62:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign Muxn_1_io_config = cfgOut[47:45]; // @[PE.scala 121:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 62:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 62:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 62:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 62:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 90:17]
  assign cfg_io_cfg_addr = io_cfg_addr[0]; // @[PE.scala 91:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 92:19]
endmodule
module GPE_49(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [3:0] alu_io_config; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 50:19]
  wire [31:0] alu_io_out; // @[PE.scala 50:19]
  wire  rf_clock; // @[PE.scala 51:18]
  wire  rf_reset; // @[PE.scala 51:18]
  wire  rf_io_en; // @[PE.scala 51:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 51:18]
  wire  DelayPipe_clock; // @[PE.scala 52:54]
  wire  DelayPipe_reset; // @[PE.scala 52:54]
  wire  DelayPipe_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 52:54]
  wire  DelayPipe_1_clock; // @[PE.scala 52:54]
  wire  DelayPipe_1_reset; // @[PE.scala 52:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 52:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 55:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 55:49]
  wire  cfg_clock; // @[PE.scala 89:19]
  wire  cfg_reset; // @[PE.scala 89:19]
  wire  cfg_io_cfg_en; // @[PE.scala 89:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 89:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 89:19]
  wire [47:0] cfg_io_out_0; // @[PE.scala 89:19]
  wire  _T_1 = 10'h89 == io_cfg_addr[11:2]; // @[PE.scala 90:48]
  wire [47:0] cfgOut = cfg_io_out_0; // @[PE.scala 96:20 PE.scala 97:10]
  ALU alu ( // @[PE.scala 50:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 51:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 52:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 52:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_16 Muxn ( // @[PE.scala 55:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_16 Muxn_1 ( // @[PE.scala 55:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_16 cfg ( // @[PE.scala 89:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 77:13]
  assign alu_io_config = cfgOut[35:32]; // @[PE.scala 100:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 71:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 71:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 75:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 76:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_io_config = cfgOut[38:36]; // @[PE.scala 113:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 70:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_1_io_config = cfgOut[41:39]; // @[PE.scala 113:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 70:23]
  assign Muxn_io_config = cfgOut[44:42]; // @[PE.scala 121:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 62:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 62:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 62:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 62:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign Muxn_1_io_config = cfgOut[47:45]; // @[PE.scala 121:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 62:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 62:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 62:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 62:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 90:17]
  assign cfg_io_cfg_addr = io_cfg_addr[0]; // @[PE.scala 91:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 92:19]
endmodule
module GPE_50(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [3:0] alu_io_config; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 50:19]
  wire [31:0] alu_io_out; // @[PE.scala 50:19]
  wire  rf_clock; // @[PE.scala 51:18]
  wire  rf_reset; // @[PE.scala 51:18]
  wire  rf_io_en; // @[PE.scala 51:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 51:18]
  wire  DelayPipe_clock; // @[PE.scala 52:54]
  wire  DelayPipe_reset; // @[PE.scala 52:54]
  wire  DelayPipe_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 52:54]
  wire  DelayPipe_1_clock; // @[PE.scala 52:54]
  wire  DelayPipe_1_reset; // @[PE.scala 52:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 52:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 55:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 55:49]
  wire  cfg_clock; // @[PE.scala 89:19]
  wire  cfg_reset; // @[PE.scala 89:19]
  wire  cfg_io_cfg_en; // @[PE.scala 89:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 89:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 89:19]
  wire [47:0] cfg_io_out_0; // @[PE.scala 89:19]
  wire  _T_1 = 10'h8a == io_cfg_addr[11:2]; // @[PE.scala 90:48]
  wire [47:0] cfgOut = cfg_io_out_0; // @[PE.scala 96:20 PE.scala 97:10]
  ALU alu ( // @[PE.scala 50:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 51:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 52:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 52:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_16 Muxn ( // @[PE.scala 55:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_16 Muxn_1 ( // @[PE.scala 55:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_16 cfg ( // @[PE.scala 89:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 77:13]
  assign alu_io_config = cfgOut[35:32]; // @[PE.scala 100:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 71:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 71:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 75:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 76:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_io_config = cfgOut[38:36]; // @[PE.scala 113:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 70:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_1_io_config = cfgOut[41:39]; // @[PE.scala 113:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 70:23]
  assign Muxn_io_config = cfgOut[44:42]; // @[PE.scala 121:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 62:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 62:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 62:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 62:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign Muxn_1_io_config = cfgOut[47:45]; // @[PE.scala 121:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 62:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 62:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 62:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 62:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 90:17]
  assign cfg_io_cfg_addr = io_cfg_addr[0]; // @[PE.scala 91:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 92:19]
endmodule
module GPE_51(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [3:0] alu_io_config; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 50:19]
  wire [31:0] alu_io_out; // @[PE.scala 50:19]
  wire  rf_clock; // @[PE.scala 51:18]
  wire  rf_reset; // @[PE.scala 51:18]
  wire  rf_io_en; // @[PE.scala 51:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 51:18]
  wire  DelayPipe_clock; // @[PE.scala 52:54]
  wire  DelayPipe_reset; // @[PE.scala 52:54]
  wire  DelayPipe_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 52:54]
  wire  DelayPipe_1_clock; // @[PE.scala 52:54]
  wire  DelayPipe_1_reset; // @[PE.scala 52:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 52:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 55:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 55:49]
  wire  cfg_clock; // @[PE.scala 89:19]
  wire  cfg_reset; // @[PE.scala 89:19]
  wire  cfg_io_cfg_en; // @[PE.scala 89:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 89:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 89:19]
  wire [47:0] cfg_io_out_0; // @[PE.scala 89:19]
  wire  _T_1 = 10'h8b == io_cfg_addr[11:2]; // @[PE.scala 90:48]
  wire [47:0] cfgOut = cfg_io_out_0; // @[PE.scala 96:20 PE.scala 97:10]
  ALU alu ( // @[PE.scala 50:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 51:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 52:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 52:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_16 Muxn ( // @[PE.scala 55:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_16 Muxn_1 ( // @[PE.scala 55:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_16 cfg ( // @[PE.scala 89:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 77:13]
  assign alu_io_config = cfgOut[35:32]; // @[PE.scala 100:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 71:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 71:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 75:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 76:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_io_config = cfgOut[38:36]; // @[PE.scala 113:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 70:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_1_io_config = cfgOut[41:39]; // @[PE.scala 113:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 70:23]
  assign Muxn_io_config = cfgOut[44:42]; // @[PE.scala 121:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 62:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 62:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 62:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 62:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign Muxn_1_io_config = cfgOut[47:45]; // @[PE.scala 121:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 62:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 62:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 62:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 62:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 90:17]
  assign cfg_io_cfg_addr = io_cfg_addr[0]; // @[PE.scala 91:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 92:19]
endmodule
module GPE_52(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [3:0] alu_io_config; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 50:19]
  wire [31:0] alu_io_out; // @[PE.scala 50:19]
  wire  rf_clock; // @[PE.scala 51:18]
  wire  rf_reset; // @[PE.scala 51:18]
  wire  rf_io_en; // @[PE.scala 51:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 51:18]
  wire  DelayPipe_clock; // @[PE.scala 52:54]
  wire  DelayPipe_reset; // @[PE.scala 52:54]
  wire  DelayPipe_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 52:54]
  wire  DelayPipe_1_clock; // @[PE.scala 52:54]
  wire  DelayPipe_1_reset; // @[PE.scala 52:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 52:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 55:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 55:49]
  wire  cfg_clock; // @[PE.scala 89:19]
  wire  cfg_reset; // @[PE.scala 89:19]
  wire  cfg_io_cfg_en; // @[PE.scala 89:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 89:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 89:19]
  wire [47:0] cfg_io_out_0; // @[PE.scala 89:19]
  wire  _T_1 = 10'h8c == io_cfg_addr[11:2]; // @[PE.scala 90:48]
  wire [47:0] cfgOut = cfg_io_out_0; // @[PE.scala 96:20 PE.scala 97:10]
  ALU alu ( // @[PE.scala 50:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 51:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 52:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 52:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_16 Muxn ( // @[PE.scala 55:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_16 Muxn_1 ( // @[PE.scala 55:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_16 cfg ( // @[PE.scala 89:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 77:13]
  assign alu_io_config = cfgOut[35:32]; // @[PE.scala 100:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 71:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 71:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 75:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 76:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_io_config = cfgOut[38:36]; // @[PE.scala 113:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 70:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_1_io_config = cfgOut[41:39]; // @[PE.scala 113:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 70:23]
  assign Muxn_io_config = cfgOut[44:42]; // @[PE.scala 121:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 62:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 62:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 62:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 62:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign Muxn_1_io_config = cfgOut[47:45]; // @[PE.scala 121:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 62:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 62:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 62:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 62:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 90:17]
  assign cfg_io_cfg_addr = io_cfg_addr[0]; // @[PE.scala 91:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 92:19]
endmodule
module GPE_53(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [3:0] alu_io_config; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 50:19]
  wire [31:0] alu_io_out; // @[PE.scala 50:19]
  wire  rf_clock; // @[PE.scala 51:18]
  wire  rf_reset; // @[PE.scala 51:18]
  wire  rf_io_en; // @[PE.scala 51:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 51:18]
  wire  DelayPipe_clock; // @[PE.scala 52:54]
  wire  DelayPipe_reset; // @[PE.scala 52:54]
  wire  DelayPipe_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 52:54]
  wire  DelayPipe_1_clock; // @[PE.scala 52:54]
  wire  DelayPipe_1_reset; // @[PE.scala 52:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 52:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 55:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 55:49]
  wire  cfg_clock; // @[PE.scala 89:19]
  wire  cfg_reset; // @[PE.scala 89:19]
  wire  cfg_io_cfg_en; // @[PE.scala 89:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 89:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 89:19]
  wire [47:0] cfg_io_out_0; // @[PE.scala 89:19]
  wire  _T_1 = 10'h8d == io_cfg_addr[11:2]; // @[PE.scala 90:48]
  wire [47:0] cfgOut = cfg_io_out_0; // @[PE.scala 96:20 PE.scala 97:10]
  ALU alu ( // @[PE.scala 50:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 51:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 52:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 52:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_16 Muxn ( // @[PE.scala 55:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_16 Muxn_1 ( // @[PE.scala 55:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_16 cfg ( // @[PE.scala 89:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 77:13]
  assign alu_io_config = cfgOut[35:32]; // @[PE.scala 100:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 71:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 71:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 75:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 76:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_io_config = cfgOut[38:36]; // @[PE.scala 113:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 70:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_1_io_config = cfgOut[41:39]; // @[PE.scala 113:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 70:23]
  assign Muxn_io_config = cfgOut[44:42]; // @[PE.scala 121:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 62:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 62:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 62:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 62:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign Muxn_1_io_config = cfgOut[47:45]; // @[PE.scala 121:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 62:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 62:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 62:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 62:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 90:17]
  assign cfg_io_cfg_addr = io_cfg_addr[0]; // @[PE.scala 91:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 92:19]
endmodule
module GPE_54(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [3:0] alu_io_config; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 50:19]
  wire [31:0] alu_io_out; // @[PE.scala 50:19]
  wire  rf_clock; // @[PE.scala 51:18]
  wire  rf_reset; // @[PE.scala 51:18]
  wire  rf_io_en; // @[PE.scala 51:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 51:18]
  wire  DelayPipe_clock; // @[PE.scala 52:54]
  wire  DelayPipe_reset; // @[PE.scala 52:54]
  wire  DelayPipe_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 52:54]
  wire  DelayPipe_1_clock; // @[PE.scala 52:54]
  wire  DelayPipe_1_reset; // @[PE.scala 52:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 52:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 55:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 55:49]
  wire  cfg_clock; // @[PE.scala 89:19]
  wire  cfg_reset; // @[PE.scala 89:19]
  wire  cfg_io_cfg_en; // @[PE.scala 89:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 89:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 89:19]
  wire [47:0] cfg_io_out_0; // @[PE.scala 89:19]
  wire  _T_1 = 10'h8e == io_cfg_addr[11:2]; // @[PE.scala 90:48]
  wire [47:0] cfgOut = cfg_io_out_0; // @[PE.scala 96:20 PE.scala 97:10]
  ALU alu ( // @[PE.scala 50:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 51:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 52:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 52:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_16 Muxn ( // @[PE.scala 55:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_16 Muxn_1 ( // @[PE.scala 55:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_16 cfg ( // @[PE.scala 89:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 77:13]
  assign alu_io_config = cfgOut[35:32]; // @[PE.scala 100:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 71:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 71:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 75:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 76:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_io_config = cfgOut[38:36]; // @[PE.scala 113:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 70:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_1_io_config = cfgOut[41:39]; // @[PE.scala 113:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 70:23]
  assign Muxn_io_config = cfgOut[44:42]; // @[PE.scala 121:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 62:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 62:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 62:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 62:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign Muxn_1_io_config = cfgOut[47:45]; // @[PE.scala 121:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 62:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 62:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 62:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 62:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 90:17]
  assign cfg_io_cfg_addr = io_cfg_addr[0]; // @[PE.scala 91:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 92:19]
endmodule
module GPE_55(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [3:0] alu_io_config; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 50:19]
  wire [31:0] alu_io_out; // @[PE.scala 50:19]
  wire  rf_clock; // @[PE.scala 51:18]
  wire  rf_reset; // @[PE.scala 51:18]
  wire  rf_io_en; // @[PE.scala 51:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 51:18]
  wire  DelayPipe_clock; // @[PE.scala 52:54]
  wire  DelayPipe_reset; // @[PE.scala 52:54]
  wire  DelayPipe_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 52:54]
  wire  DelayPipe_1_clock; // @[PE.scala 52:54]
  wire  DelayPipe_1_reset; // @[PE.scala 52:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 52:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 55:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 55:49]
  wire  cfg_clock; // @[PE.scala 89:19]
  wire  cfg_reset; // @[PE.scala 89:19]
  wire  cfg_io_cfg_en; // @[PE.scala 89:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 89:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 89:19]
  wire [47:0] cfg_io_out_0; // @[PE.scala 89:19]
  wire  _T_1 = 10'h8f == io_cfg_addr[11:2]; // @[PE.scala 90:48]
  wire [47:0] cfgOut = cfg_io_out_0; // @[PE.scala 96:20 PE.scala 97:10]
  ALU alu ( // @[PE.scala 50:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 51:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 52:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 52:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_16 Muxn ( // @[PE.scala 55:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_16 Muxn_1 ( // @[PE.scala 55:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_16 cfg ( // @[PE.scala 89:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 77:13]
  assign alu_io_config = cfgOut[35:32]; // @[PE.scala 100:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 71:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 71:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 75:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 76:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_io_config = cfgOut[38:36]; // @[PE.scala 113:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 70:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_1_io_config = cfgOut[41:39]; // @[PE.scala 113:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 70:23]
  assign Muxn_io_config = cfgOut[44:42]; // @[PE.scala 121:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 62:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 62:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 62:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 62:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign Muxn_1_io_config = cfgOut[47:45]; // @[PE.scala 121:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 62:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 62:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 62:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 62:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 90:17]
  assign cfg_io_cfg_addr = io_cfg_addr[0]; // @[PE.scala 91:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 92:19]
endmodule
module GPE_56(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [3:0] alu_io_config; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 50:19]
  wire [31:0] alu_io_out; // @[PE.scala 50:19]
  wire  rf_clock; // @[PE.scala 51:18]
  wire  rf_reset; // @[PE.scala 51:18]
  wire  rf_io_en; // @[PE.scala 51:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 51:18]
  wire  DelayPipe_clock; // @[PE.scala 52:54]
  wire  DelayPipe_reset; // @[PE.scala 52:54]
  wire  DelayPipe_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 52:54]
  wire  DelayPipe_1_clock; // @[PE.scala 52:54]
  wire  DelayPipe_1_reset; // @[PE.scala 52:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 52:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 55:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 55:49]
  wire  cfg_clock; // @[PE.scala 89:19]
  wire  cfg_reset; // @[PE.scala 89:19]
  wire  cfg_io_cfg_en; // @[PE.scala 89:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 89:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 89:19]
  wire [47:0] cfg_io_out_0; // @[PE.scala 89:19]
  wire  _T_1 = 10'h9a == io_cfg_addr[11:2]; // @[PE.scala 90:48]
  wire [47:0] cfgOut = cfg_io_out_0; // @[PE.scala 96:20 PE.scala 97:10]
  ALU alu ( // @[PE.scala 50:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 51:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 52:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 52:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_16 Muxn ( // @[PE.scala 55:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_16 Muxn_1 ( // @[PE.scala 55:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_16 cfg ( // @[PE.scala 89:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 77:13]
  assign alu_io_config = cfgOut[35:32]; // @[PE.scala 100:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 71:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 71:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 75:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 76:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_io_config = cfgOut[38:36]; // @[PE.scala 113:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 70:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_1_io_config = cfgOut[41:39]; // @[PE.scala 113:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 70:23]
  assign Muxn_io_config = cfgOut[44:42]; // @[PE.scala 121:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 62:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 62:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 62:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 62:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign Muxn_1_io_config = cfgOut[47:45]; // @[PE.scala 121:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 62:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 62:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 62:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 62:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 90:17]
  assign cfg_io_cfg_addr = io_cfg_addr[0]; // @[PE.scala 91:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 92:19]
endmodule
module GPE_57(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [3:0] alu_io_config; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 50:19]
  wire [31:0] alu_io_out; // @[PE.scala 50:19]
  wire  rf_clock; // @[PE.scala 51:18]
  wire  rf_reset; // @[PE.scala 51:18]
  wire  rf_io_en; // @[PE.scala 51:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 51:18]
  wire  DelayPipe_clock; // @[PE.scala 52:54]
  wire  DelayPipe_reset; // @[PE.scala 52:54]
  wire  DelayPipe_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 52:54]
  wire  DelayPipe_1_clock; // @[PE.scala 52:54]
  wire  DelayPipe_1_reset; // @[PE.scala 52:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 52:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 55:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 55:49]
  wire  cfg_clock; // @[PE.scala 89:19]
  wire  cfg_reset; // @[PE.scala 89:19]
  wire  cfg_io_cfg_en; // @[PE.scala 89:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 89:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 89:19]
  wire [47:0] cfg_io_out_0; // @[PE.scala 89:19]
  wire  _T_1 = 10'h9b == io_cfg_addr[11:2]; // @[PE.scala 90:48]
  wire [47:0] cfgOut = cfg_io_out_0; // @[PE.scala 96:20 PE.scala 97:10]
  ALU alu ( // @[PE.scala 50:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 51:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 52:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 52:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_16 Muxn ( // @[PE.scala 55:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_16 Muxn_1 ( // @[PE.scala 55:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_16 cfg ( // @[PE.scala 89:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 77:13]
  assign alu_io_config = cfgOut[35:32]; // @[PE.scala 100:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 71:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 71:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 75:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 76:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_io_config = cfgOut[38:36]; // @[PE.scala 113:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 70:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_1_io_config = cfgOut[41:39]; // @[PE.scala 113:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 70:23]
  assign Muxn_io_config = cfgOut[44:42]; // @[PE.scala 121:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 62:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 62:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 62:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 62:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign Muxn_1_io_config = cfgOut[47:45]; // @[PE.scala 121:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 62:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 62:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 62:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 62:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 90:17]
  assign cfg_io_cfg_addr = io_cfg_addr[0]; // @[PE.scala 91:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 92:19]
endmodule
module GPE_58(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [3:0] alu_io_config; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 50:19]
  wire [31:0] alu_io_out; // @[PE.scala 50:19]
  wire  rf_clock; // @[PE.scala 51:18]
  wire  rf_reset; // @[PE.scala 51:18]
  wire  rf_io_en; // @[PE.scala 51:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 51:18]
  wire  DelayPipe_clock; // @[PE.scala 52:54]
  wire  DelayPipe_reset; // @[PE.scala 52:54]
  wire  DelayPipe_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 52:54]
  wire  DelayPipe_1_clock; // @[PE.scala 52:54]
  wire  DelayPipe_1_reset; // @[PE.scala 52:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 52:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 55:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 55:49]
  wire  cfg_clock; // @[PE.scala 89:19]
  wire  cfg_reset; // @[PE.scala 89:19]
  wire  cfg_io_cfg_en; // @[PE.scala 89:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 89:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 89:19]
  wire [47:0] cfg_io_out_0; // @[PE.scala 89:19]
  wire  _T_1 = 10'h9c == io_cfg_addr[11:2]; // @[PE.scala 90:48]
  wire [47:0] cfgOut = cfg_io_out_0; // @[PE.scala 96:20 PE.scala 97:10]
  ALU alu ( // @[PE.scala 50:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 51:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 52:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 52:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_16 Muxn ( // @[PE.scala 55:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_16 Muxn_1 ( // @[PE.scala 55:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_16 cfg ( // @[PE.scala 89:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 77:13]
  assign alu_io_config = cfgOut[35:32]; // @[PE.scala 100:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 71:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 71:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 75:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 76:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_io_config = cfgOut[38:36]; // @[PE.scala 113:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 70:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_1_io_config = cfgOut[41:39]; // @[PE.scala 113:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 70:23]
  assign Muxn_io_config = cfgOut[44:42]; // @[PE.scala 121:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 62:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 62:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 62:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 62:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign Muxn_1_io_config = cfgOut[47:45]; // @[PE.scala 121:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 62:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 62:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 62:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 62:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 90:17]
  assign cfg_io_cfg_addr = io_cfg_addr[0]; // @[PE.scala 91:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 92:19]
endmodule
module GPE_59(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [3:0] alu_io_config; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 50:19]
  wire [31:0] alu_io_out; // @[PE.scala 50:19]
  wire  rf_clock; // @[PE.scala 51:18]
  wire  rf_reset; // @[PE.scala 51:18]
  wire  rf_io_en; // @[PE.scala 51:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 51:18]
  wire  DelayPipe_clock; // @[PE.scala 52:54]
  wire  DelayPipe_reset; // @[PE.scala 52:54]
  wire  DelayPipe_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 52:54]
  wire  DelayPipe_1_clock; // @[PE.scala 52:54]
  wire  DelayPipe_1_reset; // @[PE.scala 52:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 52:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 55:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 55:49]
  wire  cfg_clock; // @[PE.scala 89:19]
  wire  cfg_reset; // @[PE.scala 89:19]
  wire  cfg_io_cfg_en; // @[PE.scala 89:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 89:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 89:19]
  wire [47:0] cfg_io_out_0; // @[PE.scala 89:19]
  wire  _T_1 = 10'h9d == io_cfg_addr[11:2]; // @[PE.scala 90:48]
  wire [47:0] cfgOut = cfg_io_out_0; // @[PE.scala 96:20 PE.scala 97:10]
  ALU alu ( // @[PE.scala 50:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 51:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 52:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 52:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_16 Muxn ( // @[PE.scala 55:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_16 Muxn_1 ( // @[PE.scala 55:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_16 cfg ( // @[PE.scala 89:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 77:13]
  assign alu_io_config = cfgOut[35:32]; // @[PE.scala 100:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 71:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 71:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 75:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 76:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_io_config = cfgOut[38:36]; // @[PE.scala 113:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 70:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_1_io_config = cfgOut[41:39]; // @[PE.scala 113:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 70:23]
  assign Muxn_io_config = cfgOut[44:42]; // @[PE.scala 121:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 62:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 62:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 62:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 62:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign Muxn_1_io_config = cfgOut[47:45]; // @[PE.scala 121:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 62:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 62:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 62:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 62:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 90:17]
  assign cfg_io_cfg_addr = io_cfg_addr[0]; // @[PE.scala 91:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 92:19]
endmodule
module GPE_60(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [3:0] alu_io_config; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 50:19]
  wire [31:0] alu_io_out; // @[PE.scala 50:19]
  wire  rf_clock; // @[PE.scala 51:18]
  wire  rf_reset; // @[PE.scala 51:18]
  wire  rf_io_en; // @[PE.scala 51:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 51:18]
  wire  DelayPipe_clock; // @[PE.scala 52:54]
  wire  DelayPipe_reset; // @[PE.scala 52:54]
  wire  DelayPipe_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 52:54]
  wire  DelayPipe_1_clock; // @[PE.scala 52:54]
  wire  DelayPipe_1_reset; // @[PE.scala 52:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 52:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 55:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 55:49]
  wire  cfg_clock; // @[PE.scala 89:19]
  wire  cfg_reset; // @[PE.scala 89:19]
  wire  cfg_io_cfg_en; // @[PE.scala 89:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 89:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 89:19]
  wire [47:0] cfg_io_out_0; // @[PE.scala 89:19]
  wire  _T_1 = 10'h9e == io_cfg_addr[11:2]; // @[PE.scala 90:48]
  wire [47:0] cfgOut = cfg_io_out_0; // @[PE.scala 96:20 PE.scala 97:10]
  ALU alu ( // @[PE.scala 50:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 51:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 52:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 52:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_16 Muxn ( // @[PE.scala 55:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_16 Muxn_1 ( // @[PE.scala 55:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_16 cfg ( // @[PE.scala 89:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 77:13]
  assign alu_io_config = cfgOut[35:32]; // @[PE.scala 100:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 71:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 71:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 75:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 76:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_io_config = cfgOut[38:36]; // @[PE.scala 113:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 70:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_1_io_config = cfgOut[41:39]; // @[PE.scala 113:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 70:23]
  assign Muxn_io_config = cfgOut[44:42]; // @[PE.scala 121:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 62:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 62:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 62:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 62:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign Muxn_1_io_config = cfgOut[47:45]; // @[PE.scala 121:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 62:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 62:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 62:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 62:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 90:17]
  assign cfg_io_cfg_addr = io_cfg_addr[0]; // @[PE.scala 91:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 92:19]
endmodule
module GPE_61(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [3:0] alu_io_config; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 50:19]
  wire [31:0] alu_io_out; // @[PE.scala 50:19]
  wire  rf_clock; // @[PE.scala 51:18]
  wire  rf_reset; // @[PE.scala 51:18]
  wire  rf_io_en; // @[PE.scala 51:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 51:18]
  wire  DelayPipe_clock; // @[PE.scala 52:54]
  wire  DelayPipe_reset; // @[PE.scala 52:54]
  wire  DelayPipe_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 52:54]
  wire  DelayPipe_1_clock; // @[PE.scala 52:54]
  wire  DelayPipe_1_reset; // @[PE.scala 52:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 52:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 55:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 55:49]
  wire  cfg_clock; // @[PE.scala 89:19]
  wire  cfg_reset; // @[PE.scala 89:19]
  wire  cfg_io_cfg_en; // @[PE.scala 89:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 89:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 89:19]
  wire [47:0] cfg_io_out_0; // @[PE.scala 89:19]
  wire  _T_1 = 10'h9f == io_cfg_addr[11:2]; // @[PE.scala 90:48]
  wire [47:0] cfgOut = cfg_io_out_0; // @[PE.scala 96:20 PE.scala 97:10]
  ALU alu ( // @[PE.scala 50:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 51:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 52:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 52:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_16 Muxn ( // @[PE.scala 55:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_16 Muxn_1 ( // @[PE.scala 55:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_16 cfg ( // @[PE.scala 89:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 77:13]
  assign alu_io_config = cfgOut[35:32]; // @[PE.scala 100:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 71:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 71:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 75:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 76:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_io_config = cfgOut[38:36]; // @[PE.scala 113:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 70:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_1_io_config = cfgOut[41:39]; // @[PE.scala 113:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 70:23]
  assign Muxn_io_config = cfgOut[44:42]; // @[PE.scala 121:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 62:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 62:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 62:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 62:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign Muxn_1_io_config = cfgOut[47:45]; // @[PE.scala 121:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 62:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 62:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 62:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 62:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 90:17]
  assign cfg_io_cfg_addr = io_cfg_addr[0]; // @[PE.scala 91:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 92:19]
endmodule
module GPE_62(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [3:0] alu_io_config; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 50:19]
  wire [31:0] alu_io_out; // @[PE.scala 50:19]
  wire  rf_clock; // @[PE.scala 51:18]
  wire  rf_reset; // @[PE.scala 51:18]
  wire  rf_io_en; // @[PE.scala 51:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 51:18]
  wire  DelayPipe_clock; // @[PE.scala 52:54]
  wire  DelayPipe_reset; // @[PE.scala 52:54]
  wire  DelayPipe_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 52:54]
  wire  DelayPipe_1_clock; // @[PE.scala 52:54]
  wire  DelayPipe_1_reset; // @[PE.scala 52:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 52:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 55:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 55:49]
  wire  cfg_clock; // @[PE.scala 89:19]
  wire  cfg_reset; // @[PE.scala 89:19]
  wire  cfg_io_cfg_en; // @[PE.scala 89:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 89:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 89:19]
  wire [47:0] cfg_io_out_0; // @[PE.scala 89:19]
  wire  _T_1 = 10'ha0 == io_cfg_addr[11:2]; // @[PE.scala 90:48]
  wire [47:0] cfgOut = cfg_io_out_0; // @[PE.scala 96:20 PE.scala 97:10]
  ALU alu ( // @[PE.scala 50:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 51:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 52:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 52:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_16 Muxn ( // @[PE.scala 55:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_16 Muxn_1 ( // @[PE.scala 55:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_16 cfg ( // @[PE.scala 89:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 77:13]
  assign alu_io_config = cfgOut[35:32]; // @[PE.scala 100:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 71:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 71:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 75:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 76:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_io_config = cfgOut[38:36]; // @[PE.scala 113:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 70:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_1_io_config = cfgOut[41:39]; // @[PE.scala 113:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 70:23]
  assign Muxn_io_config = cfgOut[44:42]; // @[PE.scala 121:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 62:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 62:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 62:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 62:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign Muxn_1_io_config = cfgOut[47:45]; // @[PE.scala 121:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 62:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 62:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 62:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 62:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 90:17]
  assign cfg_io_cfg_addr = io_cfg_addr[0]; // @[PE.scala 91:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 92:19]
endmodule
module GPE_63(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [3:0] alu_io_config; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 50:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 50:19]
  wire [31:0] alu_io_out; // @[PE.scala 50:19]
  wire  rf_clock; // @[PE.scala 51:18]
  wire  rf_reset; // @[PE.scala 51:18]
  wire  rf_io_en; // @[PE.scala 51:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 51:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 51:18]
  wire  DelayPipe_clock; // @[PE.scala 52:54]
  wire  DelayPipe_reset; // @[PE.scala 52:54]
  wire  DelayPipe_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 52:54]
  wire  DelayPipe_1_clock; // @[PE.scala 52:54]
  wire  DelayPipe_1_reset; // @[PE.scala 52:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 52:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 52:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 52:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 55:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 55:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 55:49]
  wire  cfg_clock; // @[PE.scala 89:19]
  wire  cfg_reset; // @[PE.scala 89:19]
  wire  cfg_io_cfg_en; // @[PE.scala 89:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 89:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 89:19]
  wire [47:0] cfg_io_out_0; // @[PE.scala 89:19]
  wire  _T_1 = 10'ha1 == io_cfg_addr[11:2]; // @[PE.scala 90:48]
  wire [47:0] cfgOut = cfg_io_out_0; // @[PE.scala 96:20 PE.scala 97:10]
  ALU alu ( // @[PE.scala 50:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 51:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 52:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 52:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_16 Muxn ( // @[PE.scala 55:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_16 Muxn_1 ( // @[PE.scala 55:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_16 cfg ( // @[PE.scala 89:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 77:13]
  assign alu_io_config = cfgOut[35:32]; // @[PE.scala 100:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 71:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 71:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 75:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 76:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_io_config = cfgOut[38:36]; // @[PE.scala 113:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 70:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 69:23]
  assign DelayPipe_1_io_config = cfgOut[41:39]; // @[PE.scala 113:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 70:23]
  assign Muxn_io_config = cfgOut[44:42]; // @[PE.scala 121:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 62:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 62:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 62:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 62:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign Muxn_1_io_config = cfgOut[47:45]; // @[PE.scala 121:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 62:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 62:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 62:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 62:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 64:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 66:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 90:17]
  assign cfg_io_cfg_addr = io_cfg_addr[0]; // @[PE.scala 91:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 92:19]
endmodule
module ConfigMem_80(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [31:0] io_cfg_data,
  output [13:0] io_out_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [13:0] regs_0; // @[ConfigMem.scala 27:21]
  assign io_out_0 = regs_0; // @[ConfigMem.scala 52:45]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  regs_0 = _RAND_0[13:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      regs_0 <= 14'h0;
    end else if (io_cfg_en) begin
      regs_0 <= io_cfg_data[13:0];
    end
  end
endmodule
module Muxn_145(
  input  [1:0]  io_config,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  output [31:0] io_out
);
  wire  _T_2 = 2'h1 == io_config; // @[Mux.scala 80:60]
  wire [31:0] _T_3 = _T_2 ? io_in_1 : io_in_0; // @[Mux.scala 80:57]
  wire  _T_4 = 2'h2 == io_config; // @[Mux.scala 80:60]
  assign io_out = _T_4 ? io_in_2 : _T_3; // @[Multiplexer.scala 20:10]
endmodule
module Muxn_147(
  input  [2:0]  io_config,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  output [31:0] io_out
);
  wire  _T_2 = 3'h1 == io_config; // @[Mux.scala 80:60]
  wire [31:0] _T_3 = _T_2 ? io_in_1 : io_in_0; // @[Mux.scala 80:57]
  wire  _T_4 = 3'h2 == io_config; // @[Mux.scala 80:60]
  wire [31:0] _T_5 = _T_4 ? io_in_2 : _T_3; // @[Mux.scala 80:57]
  wire  _T_6 = 3'h3 == io_config; // @[Mux.scala 80:60]
  wire [31:0] _T_7 = _T_6 ? io_in_3 : _T_5; // @[Mux.scala 80:57]
  wire  _T_8 = 3'h4 == io_config; // @[Mux.scala 80:60]
  assign io_out = _T_8 ? io_in_4 : _T_7; // @[Multiplexer.scala 20:10]
endmodule
module Muxn_148(
  input  [1:0]  io_config,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  output [31:0] io_out
);
  wire  _T = 2'h1 == io_config; // @[Mux.scala 80:60]
  wire [31:0] _T_1 = _T ? io_in_1 : io_in_0; // @[Mux.scala 80:57]
  wire  _T_2 = 2'h2 == io_config; // @[Mux.scala 80:60]
  wire [31:0] _T_3 = _T_2 ? io_in_2 : _T_1; // @[Mux.scala 80:57]
  wire  _T_4 = 2'h3 == io_config; // @[Mux.scala 80:60]
  assign io_out = _T_4 ? io_in_3 : _T_3; // @[Multiplexer.scala 20:10]
endmodule
module GIB(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNE_0,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
  wire  ConfigMem_clock; // @[Interconnect.scala 463:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 463:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 463:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 463:21]
  wire [13:0] ConfigMem_io_out_0; // @[Interconnect.scala 463:21]
  wire  Muxn_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_3_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_6_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 473:25]
  wire  _T_1 = 10'h13 == io_cfg_addr[11:2]; // @[Interconnect.scala 464:50]
  ConfigMem_80 ConfigMem ( // @[Interconnect.scala 463:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn Muxn ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_out(Muxn_io_out)
  );
  Muxn_145 Muxn_1 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_out(Muxn_1_io_out)
  );
  Muxn_145 Muxn_2 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_out(Muxn_2_io_out)
  );
  Muxn_147 Muxn_3 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_in_3(Muxn_3_io_in_3),
    .io_in_4(Muxn_3_io_in_4),
    .io_out(Muxn_3_io_out)
  );
  Muxn_148 Muxn_4 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_in_3(Muxn_4_io_in_3),
    .io_out(Muxn_4_io_out)
  );
  Muxn_145 Muxn_5 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_out(Muxn_5_io_out)
  );
  Muxn_148 Muxn_6 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_out(Muxn_6_io_out)
  );
  assign io_ipinNE_0 = Muxn_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinSE_0 = Muxn_1_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSE_1 = Muxn_2_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_otrackE_0 = Muxn_5_io_out; // @[Interconnect.scala 432:21 Interconnect.scala 479:45]
  assign io_otrackS_0 = Muxn_6_io_out; // @[Interconnect.scala 433:21 Interconnect.scala 479:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 464:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 466:21]
  assign Muxn_io_config = ConfigMem_io_out_0[0]; // @[Interconnect.scala 483:23]
  assign Muxn_io_in_0 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_1 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[2:1]; // @[Interconnect.scala 483:23]
  assign Muxn_1_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_1 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_2 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[4:3]; // @[Interconnect.scala 483:23]
  assign Muxn_2_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_1 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_2 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:5]; // @[Interconnect.scala 483:23]
  assign Muxn_3_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_2 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 483:23]
  assign Muxn_4_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_1 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 483:23]
  assign Muxn_5_io_in_0 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_1 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_2 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[13:12]; // @[Interconnect.scala 483:23]
  assign Muxn_6_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_1 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_2 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
endmodule
module ConfigMem_81(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [31:0] io_cfg_data,
  output [23:0] io_out_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [23:0] regs_0; // @[ConfigMem.scala 27:21]
  assign io_out_0 = regs_0; // @[ConfigMem.scala 52:45]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  regs_0 = _RAND_0[23:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      regs_0 <= 24'h0;
    end else if (io_cfg_en) begin
      regs_0 <= io_cfg_data[23:0];
    end
  end
endmodule
module GIB_1(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire  ConfigMem_clock; // @[Interconnect.scala 463:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 463:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 463:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 463:21]
  wire [23:0] ConfigMem_io_out_0; // @[Interconnect.scala 463:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_6_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_7_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 473:25]
  wire  _T_1 = 10'h14 == io_cfg_addr[11:2]; // @[Interconnect.scala 464:50]
  reg [31:0] _T_10; // @[Interconnect.scala 477:55]
  reg [31:0] _T_14; // @[Interconnect.scala 477:55]
  reg [31:0] _T_16; // @[Interconnect.scala 477:55]
  ConfigMem_81 ConfigMem ( // @[Interconnect.scala 463:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_148 Muxn ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_out(Muxn_io_out)
  );
  Muxn_148 Muxn_1 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_out(Muxn_1_io_out)
  );
  Muxn_148 Muxn_2 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_in_3(Muxn_2_io_in_3),
    .io_out(Muxn_2_io_out)
  );
  Muxn_148 Muxn_3 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_in_3(Muxn_3_io_in_3),
    .io_out(Muxn_3_io_out)
  );
  Muxn_148 Muxn_4 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_in_3(Muxn_4_io_in_3),
    .io_out(Muxn_4_io_out)
  );
  Muxn_148 Muxn_5 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_in_3(Muxn_5_io_in_3),
    .io_out(Muxn_5_io_out)
  );
  Muxn_147 Muxn_6 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_in_4(Muxn_6_io_in_4),
    .io_out(Muxn_6_io_out)
  );
  Muxn_147 Muxn_7 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_in_4(Muxn_7_io_in_4),
    .io_out(Muxn_7_io_out)
  );
  Muxn_147 Muxn_8 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_147 Muxn_9 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNE_0 = Muxn_1_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinSE_0 = Muxn_2_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSE_1 = Muxn_3_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSW_0 = Muxn_4_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_ipinSW_1 = Muxn_5_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_otrackW_0 = _T_10; // @[Interconnect.scala 430:21 Interconnect.scala 477:45]
  assign io_otrackE_0 = _T_14; // @[Interconnect.scala 432:21 Interconnect.scala 477:45]
  assign io_otrackS_0 = _T_16; // @[Interconnect.scala 433:21 Interconnect.scala 477:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 464:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 466:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 483:23]
  assign Muxn_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 483:23]
  assign Muxn_1_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 483:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_3 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 483:23]
  assign Muxn_3_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_3 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 483:23]
  assign Muxn_4_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_2 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 483:23]
  assign Muxn_5_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_2 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[14:12]; // @[Interconnect.scala 483:23]
  assign Muxn_6_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_2 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[17:15]; // @[Interconnect.scala 483:23]
  assign Muxn_7_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[20:18]; // @[Interconnect.scala 483:23]
  assign Muxn_8_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_3 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[23:21]; // @[Interconnect.scala 483:23]
  assign Muxn_9_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_3 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_4 = io_itrackE_0; // @[Interconnect.scala 475:63]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_10 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  _T_14 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  _T_16 = _RAND_2[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_10 <= Muxn_6_io_out;
    _T_14 <= Muxn_8_io_out;
    _T_16 <= Muxn_9_io_out;
  end
endmodule
module GIB_2(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
  wire  ConfigMem_clock; // @[Interconnect.scala 463:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 463:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 463:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 463:21]
  wire [23:0] ConfigMem_io_out_0; // @[Interconnect.scala 463:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_6_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_7_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 473:25]
  wire  _T_1 = 10'h15 == io_cfg_addr[11:2]; // @[Interconnect.scala 464:50]
  ConfigMem_81 ConfigMem ( // @[Interconnect.scala 463:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_148 Muxn ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_out(Muxn_io_out)
  );
  Muxn_148 Muxn_1 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_out(Muxn_1_io_out)
  );
  Muxn_148 Muxn_2 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_in_3(Muxn_2_io_in_3),
    .io_out(Muxn_2_io_out)
  );
  Muxn_148 Muxn_3 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_in_3(Muxn_3_io_in_3),
    .io_out(Muxn_3_io_out)
  );
  Muxn_148 Muxn_4 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_in_3(Muxn_4_io_in_3),
    .io_out(Muxn_4_io_out)
  );
  Muxn_148 Muxn_5 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_in_3(Muxn_5_io_in_3),
    .io_out(Muxn_5_io_out)
  );
  Muxn_147 Muxn_6 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_in_4(Muxn_6_io_in_4),
    .io_out(Muxn_6_io_out)
  );
  Muxn_147 Muxn_7 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_in_4(Muxn_7_io_in_4),
    .io_out(Muxn_7_io_out)
  );
  Muxn_147 Muxn_8 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_147 Muxn_9 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNE_0 = Muxn_1_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinSE_0 = Muxn_2_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSE_1 = Muxn_3_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSW_0 = Muxn_4_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_ipinSW_1 = Muxn_5_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_otrackW_0 = Muxn_6_io_out; // @[Interconnect.scala 430:21 Interconnect.scala 479:45]
  assign io_otrackE_0 = Muxn_8_io_out; // @[Interconnect.scala 432:21 Interconnect.scala 479:45]
  assign io_otrackS_0 = Muxn_9_io_out; // @[Interconnect.scala 433:21 Interconnect.scala 479:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 464:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 466:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 483:23]
  assign Muxn_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 483:23]
  assign Muxn_1_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 483:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_3 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 483:23]
  assign Muxn_3_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_3 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 483:23]
  assign Muxn_4_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_2 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 483:23]
  assign Muxn_5_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_2 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[14:12]; // @[Interconnect.scala 483:23]
  assign Muxn_6_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_2 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[17:15]; // @[Interconnect.scala 483:23]
  assign Muxn_7_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[20:18]; // @[Interconnect.scala 483:23]
  assign Muxn_8_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_3 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[23:21]; // @[Interconnect.scala 483:23]
  assign Muxn_9_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_3 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_4 = io_itrackE_0; // @[Interconnect.scala 475:63]
endmodule
module GIB_3(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire  ConfigMem_clock; // @[Interconnect.scala 463:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 463:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 463:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 463:21]
  wire [23:0] ConfigMem_io_out_0; // @[Interconnect.scala 463:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_6_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_7_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 473:25]
  wire  _T_1 = 10'h16 == io_cfg_addr[11:2]; // @[Interconnect.scala 464:50]
  reg [31:0] _T_10; // @[Interconnect.scala 477:55]
  reg [31:0] _T_14; // @[Interconnect.scala 477:55]
  reg [31:0] _T_16; // @[Interconnect.scala 477:55]
  ConfigMem_81 ConfigMem ( // @[Interconnect.scala 463:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_148 Muxn ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_out(Muxn_io_out)
  );
  Muxn_148 Muxn_1 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_out(Muxn_1_io_out)
  );
  Muxn_148 Muxn_2 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_in_3(Muxn_2_io_in_3),
    .io_out(Muxn_2_io_out)
  );
  Muxn_148 Muxn_3 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_in_3(Muxn_3_io_in_3),
    .io_out(Muxn_3_io_out)
  );
  Muxn_148 Muxn_4 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_in_3(Muxn_4_io_in_3),
    .io_out(Muxn_4_io_out)
  );
  Muxn_148 Muxn_5 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_in_3(Muxn_5_io_in_3),
    .io_out(Muxn_5_io_out)
  );
  Muxn_147 Muxn_6 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_in_4(Muxn_6_io_in_4),
    .io_out(Muxn_6_io_out)
  );
  Muxn_147 Muxn_7 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_in_4(Muxn_7_io_in_4),
    .io_out(Muxn_7_io_out)
  );
  Muxn_147 Muxn_8 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_147 Muxn_9 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNE_0 = Muxn_1_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinSE_0 = Muxn_2_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSE_1 = Muxn_3_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSW_0 = Muxn_4_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_ipinSW_1 = Muxn_5_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_otrackW_0 = _T_10; // @[Interconnect.scala 430:21 Interconnect.scala 477:45]
  assign io_otrackE_0 = _T_14; // @[Interconnect.scala 432:21 Interconnect.scala 477:45]
  assign io_otrackS_0 = _T_16; // @[Interconnect.scala 433:21 Interconnect.scala 477:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 464:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 466:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 483:23]
  assign Muxn_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 483:23]
  assign Muxn_1_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 483:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_3 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 483:23]
  assign Muxn_3_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_3 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 483:23]
  assign Muxn_4_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_2 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 483:23]
  assign Muxn_5_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_2 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[14:12]; // @[Interconnect.scala 483:23]
  assign Muxn_6_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_2 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[17:15]; // @[Interconnect.scala 483:23]
  assign Muxn_7_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[20:18]; // @[Interconnect.scala 483:23]
  assign Muxn_8_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_3 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[23:21]; // @[Interconnect.scala 483:23]
  assign Muxn_9_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_3 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_4 = io_itrackE_0; // @[Interconnect.scala 475:63]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_10 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  _T_14 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  _T_16 = _RAND_2[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_10 <= Muxn_6_io_out;
    _T_14 <= Muxn_8_io_out;
    _T_16 <= Muxn_9_io_out;
  end
endmodule
module GIB_4(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
  wire  ConfigMem_clock; // @[Interconnect.scala 463:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 463:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 463:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 463:21]
  wire [23:0] ConfigMem_io_out_0; // @[Interconnect.scala 463:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_6_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_7_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 473:25]
  wire  _T_1 = 10'h17 == io_cfg_addr[11:2]; // @[Interconnect.scala 464:50]
  ConfigMem_81 ConfigMem ( // @[Interconnect.scala 463:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_148 Muxn ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_out(Muxn_io_out)
  );
  Muxn_148 Muxn_1 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_out(Muxn_1_io_out)
  );
  Muxn_148 Muxn_2 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_in_3(Muxn_2_io_in_3),
    .io_out(Muxn_2_io_out)
  );
  Muxn_148 Muxn_3 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_in_3(Muxn_3_io_in_3),
    .io_out(Muxn_3_io_out)
  );
  Muxn_148 Muxn_4 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_in_3(Muxn_4_io_in_3),
    .io_out(Muxn_4_io_out)
  );
  Muxn_148 Muxn_5 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_in_3(Muxn_5_io_in_3),
    .io_out(Muxn_5_io_out)
  );
  Muxn_147 Muxn_6 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_in_4(Muxn_6_io_in_4),
    .io_out(Muxn_6_io_out)
  );
  Muxn_147 Muxn_7 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_in_4(Muxn_7_io_in_4),
    .io_out(Muxn_7_io_out)
  );
  Muxn_147 Muxn_8 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_147 Muxn_9 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNE_0 = Muxn_1_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinSE_0 = Muxn_2_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSE_1 = Muxn_3_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSW_0 = Muxn_4_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_ipinSW_1 = Muxn_5_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_otrackW_0 = Muxn_6_io_out; // @[Interconnect.scala 430:21 Interconnect.scala 479:45]
  assign io_otrackE_0 = Muxn_8_io_out; // @[Interconnect.scala 432:21 Interconnect.scala 479:45]
  assign io_otrackS_0 = Muxn_9_io_out; // @[Interconnect.scala 433:21 Interconnect.scala 479:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 464:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 466:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 483:23]
  assign Muxn_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 483:23]
  assign Muxn_1_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 483:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_3 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 483:23]
  assign Muxn_3_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_3 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 483:23]
  assign Muxn_4_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_2 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 483:23]
  assign Muxn_5_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_2 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[14:12]; // @[Interconnect.scala 483:23]
  assign Muxn_6_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_2 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[17:15]; // @[Interconnect.scala 483:23]
  assign Muxn_7_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[20:18]; // @[Interconnect.scala 483:23]
  assign Muxn_8_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_3 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[23:21]; // @[Interconnect.scala 483:23]
  assign Muxn_9_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_3 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_4 = io_itrackE_0; // @[Interconnect.scala 475:63]
endmodule
module GIB_5(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire  ConfigMem_clock; // @[Interconnect.scala 463:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 463:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 463:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 463:21]
  wire [23:0] ConfigMem_io_out_0; // @[Interconnect.scala 463:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_6_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_7_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 473:25]
  wire  _T_1 = 10'h18 == io_cfg_addr[11:2]; // @[Interconnect.scala 464:50]
  reg [31:0] _T_10; // @[Interconnect.scala 477:55]
  reg [31:0] _T_14; // @[Interconnect.scala 477:55]
  reg [31:0] _T_16; // @[Interconnect.scala 477:55]
  ConfigMem_81 ConfigMem ( // @[Interconnect.scala 463:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_148 Muxn ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_out(Muxn_io_out)
  );
  Muxn_148 Muxn_1 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_out(Muxn_1_io_out)
  );
  Muxn_148 Muxn_2 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_in_3(Muxn_2_io_in_3),
    .io_out(Muxn_2_io_out)
  );
  Muxn_148 Muxn_3 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_in_3(Muxn_3_io_in_3),
    .io_out(Muxn_3_io_out)
  );
  Muxn_148 Muxn_4 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_in_3(Muxn_4_io_in_3),
    .io_out(Muxn_4_io_out)
  );
  Muxn_148 Muxn_5 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_in_3(Muxn_5_io_in_3),
    .io_out(Muxn_5_io_out)
  );
  Muxn_147 Muxn_6 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_in_4(Muxn_6_io_in_4),
    .io_out(Muxn_6_io_out)
  );
  Muxn_147 Muxn_7 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_in_4(Muxn_7_io_in_4),
    .io_out(Muxn_7_io_out)
  );
  Muxn_147 Muxn_8 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_147 Muxn_9 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNE_0 = Muxn_1_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinSE_0 = Muxn_2_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSE_1 = Muxn_3_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSW_0 = Muxn_4_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_ipinSW_1 = Muxn_5_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_otrackW_0 = _T_10; // @[Interconnect.scala 430:21 Interconnect.scala 477:45]
  assign io_otrackE_0 = _T_14; // @[Interconnect.scala 432:21 Interconnect.scala 477:45]
  assign io_otrackS_0 = _T_16; // @[Interconnect.scala 433:21 Interconnect.scala 477:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 464:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 466:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 483:23]
  assign Muxn_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 483:23]
  assign Muxn_1_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 483:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_3 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 483:23]
  assign Muxn_3_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_3 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 483:23]
  assign Muxn_4_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_2 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 483:23]
  assign Muxn_5_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_2 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[14:12]; // @[Interconnect.scala 483:23]
  assign Muxn_6_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_2 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[17:15]; // @[Interconnect.scala 483:23]
  assign Muxn_7_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[20:18]; // @[Interconnect.scala 483:23]
  assign Muxn_8_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_3 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[23:21]; // @[Interconnect.scala 483:23]
  assign Muxn_9_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_3 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_4 = io_itrackE_0; // @[Interconnect.scala 475:63]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_10 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  _T_14 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  _T_16 = _RAND_2[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_10 <= Muxn_6_io_out;
    _T_14 <= Muxn_8_io_out;
    _T_16 <= Muxn_9_io_out;
  end
endmodule
module GIB_6(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
  wire  ConfigMem_clock; // @[Interconnect.scala 463:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 463:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 463:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 463:21]
  wire [23:0] ConfigMem_io_out_0; // @[Interconnect.scala 463:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_6_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_7_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 473:25]
  wire  _T_1 = 10'h19 == io_cfg_addr[11:2]; // @[Interconnect.scala 464:50]
  ConfigMem_81 ConfigMem ( // @[Interconnect.scala 463:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_148 Muxn ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_out(Muxn_io_out)
  );
  Muxn_148 Muxn_1 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_out(Muxn_1_io_out)
  );
  Muxn_148 Muxn_2 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_in_3(Muxn_2_io_in_3),
    .io_out(Muxn_2_io_out)
  );
  Muxn_148 Muxn_3 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_in_3(Muxn_3_io_in_3),
    .io_out(Muxn_3_io_out)
  );
  Muxn_148 Muxn_4 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_in_3(Muxn_4_io_in_3),
    .io_out(Muxn_4_io_out)
  );
  Muxn_148 Muxn_5 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_in_3(Muxn_5_io_in_3),
    .io_out(Muxn_5_io_out)
  );
  Muxn_147 Muxn_6 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_in_4(Muxn_6_io_in_4),
    .io_out(Muxn_6_io_out)
  );
  Muxn_147 Muxn_7 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_in_4(Muxn_7_io_in_4),
    .io_out(Muxn_7_io_out)
  );
  Muxn_147 Muxn_8 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_147 Muxn_9 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNE_0 = Muxn_1_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinSE_0 = Muxn_2_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSE_1 = Muxn_3_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSW_0 = Muxn_4_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_ipinSW_1 = Muxn_5_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_otrackW_0 = Muxn_6_io_out; // @[Interconnect.scala 430:21 Interconnect.scala 479:45]
  assign io_otrackE_0 = Muxn_8_io_out; // @[Interconnect.scala 432:21 Interconnect.scala 479:45]
  assign io_otrackS_0 = Muxn_9_io_out; // @[Interconnect.scala 433:21 Interconnect.scala 479:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 464:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 466:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 483:23]
  assign Muxn_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 483:23]
  assign Muxn_1_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 483:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_3 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 483:23]
  assign Muxn_3_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_3 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 483:23]
  assign Muxn_4_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_2 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 483:23]
  assign Muxn_5_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_2 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[14:12]; // @[Interconnect.scala 483:23]
  assign Muxn_6_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_2 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[17:15]; // @[Interconnect.scala 483:23]
  assign Muxn_7_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[20:18]; // @[Interconnect.scala 483:23]
  assign Muxn_8_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_3 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[23:21]; // @[Interconnect.scala 483:23]
  assign Muxn_9_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_3 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_4 = io_itrackE_0; // @[Interconnect.scala 475:63]
endmodule
module GIB_7(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire  ConfigMem_clock; // @[Interconnect.scala 463:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 463:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 463:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 463:21]
  wire [23:0] ConfigMem_io_out_0; // @[Interconnect.scala 463:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_6_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_7_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 473:25]
  wire  _T_1 = 10'h1a == io_cfg_addr[11:2]; // @[Interconnect.scala 464:50]
  reg [31:0] _T_10; // @[Interconnect.scala 477:55]
  reg [31:0] _T_14; // @[Interconnect.scala 477:55]
  reg [31:0] _T_16; // @[Interconnect.scala 477:55]
  ConfigMem_81 ConfigMem ( // @[Interconnect.scala 463:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_148 Muxn ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_out(Muxn_io_out)
  );
  Muxn_148 Muxn_1 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_out(Muxn_1_io_out)
  );
  Muxn_148 Muxn_2 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_in_3(Muxn_2_io_in_3),
    .io_out(Muxn_2_io_out)
  );
  Muxn_148 Muxn_3 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_in_3(Muxn_3_io_in_3),
    .io_out(Muxn_3_io_out)
  );
  Muxn_148 Muxn_4 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_in_3(Muxn_4_io_in_3),
    .io_out(Muxn_4_io_out)
  );
  Muxn_148 Muxn_5 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_in_3(Muxn_5_io_in_3),
    .io_out(Muxn_5_io_out)
  );
  Muxn_147 Muxn_6 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_in_4(Muxn_6_io_in_4),
    .io_out(Muxn_6_io_out)
  );
  Muxn_147 Muxn_7 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_in_4(Muxn_7_io_in_4),
    .io_out(Muxn_7_io_out)
  );
  Muxn_147 Muxn_8 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_147 Muxn_9 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNE_0 = Muxn_1_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinSE_0 = Muxn_2_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSE_1 = Muxn_3_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSW_0 = Muxn_4_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_ipinSW_1 = Muxn_5_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_otrackW_0 = _T_10; // @[Interconnect.scala 430:21 Interconnect.scala 477:45]
  assign io_otrackE_0 = _T_14; // @[Interconnect.scala 432:21 Interconnect.scala 477:45]
  assign io_otrackS_0 = _T_16; // @[Interconnect.scala 433:21 Interconnect.scala 477:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 464:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 466:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 483:23]
  assign Muxn_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 483:23]
  assign Muxn_1_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 483:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_3 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 483:23]
  assign Muxn_3_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_3 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 483:23]
  assign Muxn_4_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_2 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 483:23]
  assign Muxn_5_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_2 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[14:12]; // @[Interconnect.scala 483:23]
  assign Muxn_6_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_2 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[17:15]; // @[Interconnect.scala 483:23]
  assign Muxn_7_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[20:18]; // @[Interconnect.scala 483:23]
  assign Muxn_8_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_3 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[23:21]; // @[Interconnect.scala 483:23]
  assign Muxn_9_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_3 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_4 = io_itrackE_0; // @[Interconnect.scala 475:63]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_10 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  _T_14 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  _T_16 = _RAND_2[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_10 <= Muxn_6_io_out;
    _T_14 <= Muxn_8_io_out;
    _T_16 <= Muxn_9_io_out;
  end
endmodule
module ConfigMem_88(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [31:0] io_cfg_data,
  output [12:0] io_out_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [12:0] regs_0; // @[ConfigMem.scala 27:21]
  assign io_out_0 = regs_0; // @[ConfigMem.scala 52:45]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  regs_0 = _RAND_0[12:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      regs_0 <= 13'h0;
    end else if (io_cfg_en) begin
      regs_0 <= io_cfg_data[12:0];
    end
  end
endmodule
module GIB_8(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
  wire  ConfigMem_clock; // @[Interconnect.scala 463:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 463:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 463:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 463:21]
  wire [12:0] ConfigMem_io_out_0; // @[Interconnect.scala 463:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 473:25]
  wire  Muxn_1_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 473:25]
  wire  Muxn_2_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_5_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_6_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 473:25]
  wire  _T_1 = 10'h1b == io_cfg_addr[11:2]; // @[Interconnect.scala 464:50]
  ConfigMem_88 ConfigMem ( // @[Interconnect.scala 463:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_145 Muxn ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_out(Muxn_io_out)
  );
  Muxn Muxn_1 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_out(Muxn_1_io_out)
  );
  Muxn Muxn_2 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_out(Muxn_2_io_out)
  );
  Muxn_145 Muxn_3 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_out(Muxn_3_io_out)
  );
  Muxn_148 Muxn_4 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_in_3(Muxn_4_io_in_3),
    .io_out(Muxn_4_io_out)
  );
  Muxn_147 Muxn_5 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_in_3(Muxn_5_io_in_3),
    .io_in_4(Muxn_5_io_in_4),
    .io_out(Muxn_5_io_out)
  );
  Muxn_148 Muxn_6 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_out(Muxn_6_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinSW_0 = Muxn_1_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_ipinSW_1 = Muxn_2_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_otrackW_0 = Muxn_3_io_out; // @[Interconnect.scala 430:21 Interconnect.scala 479:45]
  assign io_otrackS_0 = Muxn_6_io_out; // @[Interconnect.scala 433:21 Interconnect.scala 479:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 464:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 466:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 483:23]
  assign Muxn_io_in_0 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_1 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_2 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[2]; // @[Interconnect.scala 483:23]
  assign Muxn_1_io_in_0 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_1 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[3]; // @[Interconnect.scala 483:23]
  assign Muxn_2_io_in_0 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_1 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 483:23]
  assign Muxn_3_io_in_0 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_1 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_2 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 483:23]
  assign Muxn_4_io_in_0 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_1 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_2 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[10:8]; // @[Interconnect.scala 483:23]
  assign Muxn_5_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_3 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[12:11]; // @[Interconnect.scala 483:23]
  assign Muxn_6_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_1 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_2 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_3 = 32'h0; // @[Interconnect.scala 475:63]
endmodule
module ConfigMem_89(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [31:0] io_cfg_data,
  output [14:0] io_out_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [14:0] regs_0; // @[ConfigMem.scala 27:21]
  assign io_out_0 = regs_0; // @[ConfigMem.scala 52:45]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  regs_0 = _RAND_0[14:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      regs_0 <= 15'h0;
    end else if (io_cfg_en) begin
      regs_0 <= io_cfg_data[14:0];
    end
  end
endmodule
module GIB_9(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire  ConfigMem_clock; // @[Interconnect.scala 463:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 463:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 463:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 463:21]
  wire [14:0] ConfigMem_io_out_0; // @[Interconnect.scala 463:21]
  wire  Muxn_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 473:25]
  wire  Muxn_1_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_4_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_6_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_7_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 473:25]
  wire  _T_1 = 10'h25 == io_cfg_addr[11:2]; // @[Interconnect.scala 464:50]
  reg [31:0] _T_10; // @[Interconnect.scala 477:55]
  reg [31:0] _T_12; // @[Interconnect.scala 477:55]
  reg [31:0] _T_14; // @[Interconnect.scala 477:55]
  ConfigMem_89 ConfigMem ( // @[Interconnect.scala 463:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn Muxn ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_out(Muxn_io_out)
  );
  Muxn Muxn_1 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_out(Muxn_1_io_out)
  );
  Muxn_145 Muxn_2 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_out(Muxn_2_io_out)
  );
  Muxn_145 Muxn_3 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_out(Muxn_3_io_out)
  );
  Muxn_147 Muxn_4 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_in_3(Muxn_4_io_in_3),
    .io_in_4(Muxn_4_io_in_4),
    .io_out(Muxn_4_io_out)
  );
  Muxn_148 Muxn_5 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_in_3(Muxn_5_io_in_3),
    .io_out(Muxn_5_io_out)
  );
  Muxn_145 Muxn_6 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_out(Muxn_6_io_out)
  );
  Muxn_148 Muxn_7 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_out(Muxn_7_io_out)
  );
  assign io_ipinNE_0 = Muxn_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinNE_1 = Muxn_1_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinSE_0 = Muxn_2_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSE_1 = Muxn_3_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_otrackN_0 = _T_10; // @[Interconnect.scala 431:21 Interconnect.scala 477:45]
  assign io_otrackE_0 = _T_12; // @[Interconnect.scala 432:21 Interconnect.scala 477:45]
  assign io_otrackS_0 = _T_14; // @[Interconnect.scala 433:21 Interconnect.scala 477:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 464:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 466:21]
  assign Muxn_io_config = ConfigMem_io_out_0[0]; // @[Interconnect.scala 483:23]
  assign Muxn_io_in_0 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_1 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[1]; // @[Interconnect.scala 483:23]
  assign Muxn_1_io_in_0 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_1 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 483:23]
  assign Muxn_2_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_1 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 483:23]
  assign Muxn_3_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_1 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[8:6]; // @[Interconnect.scala 483:23]
  assign Muxn_4_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[10:9]; // @[Interconnect.scala 483:23]
  assign Muxn_5_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_1 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[12:11]; // @[Interconnect.scala 483:23]
  assign Muxn_6_io_in_0 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_1 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_2 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[14:13]; // @[Interconnect.scala 483:23]
  assign Muxn_7_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_1 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_10 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  _T_12 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  _T_14 = _RAND_2[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_10 <= Muxn_5_io_out;
    _T_12 <= Muxn_6_io_out;
    _T_14 <= Muxn_7_io_out;
  end
endmodule
module ConfigMem_90(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [31:0] io_cfg_data,
  output [27:0] io_out_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [27:0] regs_0; // @[ConfigMem.scala 27:21]
  assign io_out_0 = regs_0; // @[ConfigMem.scala 52:45]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  regs_0 = _RAND_0[27:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      regs_0 <= 28'h0;
    end else if (io_cfg_en) begin
      regs_0 <= io_cfg_data[27:0];
    end
  end
endmodule
module GIB_10(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
  wire  ConfigMem_clock; // @[Interconnect.scala 463:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 463:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 463:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 463:21]
  wire [27:0] ConfigMem_io_out_0; // @[Interconnect.scala 463:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_6_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_7_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_10_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_11_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_out; // @[Interconnect.scala 473:25]
  wire  _T_1 = 10'h26 == io_cfg_addr[11:2]; // @[Interconnect.scala 464:50]
  ConfigMem_90 ConfigMem ( // @[Interconnect.scala 463:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_148 Muxn ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_out(Muxn_io_out)
  );
  Muxn_148 Muxn_1 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_out(Muxn_1_io_out)
  );
  Muxn_148 Muxn_2 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_in_3(Muxn_2_io_in_3),
    .io_out(Muxn_2_io_out)
  );
  Muxn_148 Muxn_3 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_in_3(Muxn_3_io_in_3),
    .io_out(Muxn_3_io_out)
  );
  Muxn_148 Muxn_4 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_in_3(Muxn_4_io_in_3),
    .io_out(Muxn_4_io_out)
  );
  Muxn_148 Muxn_5 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_in_3(Muxn_5_io_in_3),
    .io_out(Muxn_5_io_out)
  );
  Muxn_148 Muxn_6 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_out(Muxn_6_io_out)
  );
  Muxn_148 Muxn_7 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_out(Muxn_7_io_out)
  );
  Muxn_147 Muxn_8 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_147 Muxn_9 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  Muxn_147 Muxn_10 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_10_io_config),
    .io_in_0(Muxn_10_io_in_0),
    .io_in_1(Muxn_10_io_in_1),
    .io_in_2(Muxn_10_io_in_2),
    .io_in_3(Muxn_10_io_in_3),
    .io_in_4(Muxn_10_io_in_4),
    .io_out(Muxn_10_io_out)
  );
  Muxn_147 Muxn_11 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_11_io_config),
    .io_in_0(Muxn_11_io_in_0),
    .io_in_1(Muxn_11_io_in_1),
    .io_in_2(Muxn_11_io_in_2),
    .io_in_3(Muxn_11_io_in_3),
    .io_in_4(Muxn_11_io_in_4),
    .io_out(Muxn_11_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNE_0 = Muxn_2_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinNE_1 = Muxn_3_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinSE_0 = Muxn_4_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSE_1 = Muxn_5_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSW_0 = Muxn_6_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_ipinSW_1 = Muxn_7_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_otrackW_0 = Muxn_8_io_out; // @[Interconnect.scala 430:21 Interconnect.scala 479:45]
  assign io_otrackN_0 = Muxn_9_io_out; // @[Interconnect.scala 431:21 Interconnect.scala 479:45]
  assign io_otrackE_0 = Muxn_10_io_out; // @[Interconnect.scala 432:21 Interconnect.scala 479:45]
  assign io_otrackS_0 = Muxn_11_io_out; // @[Interconnect.scala 433:21 Interconnect.scala 479:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 464:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 466:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 483:23]
  assign Muxn_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 483:23]
  assign Muxn_1_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 483:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 483:23]
  assign Muxn_3_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 483:23]
  assign Muxn_4_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 483:23]
  assign Muxn_5_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[13:12]; // @[Interconnect.scala 483:23]
  assign Muxn_6_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[15:14]; // @[Interconnect.scala 483:23]
  assign Muxn_7_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[18:16]; // @[Interconnect.scala 483:23]
  assign Muxn_8_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[21:19]; // @[Interconnect.scala 483:23]
  assign Muxn_9_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_config = ConfigMem_io_out_0[24:22]; // @[Interconnect.scala 483:23]
  assign Muxn_10_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_config = ConfigMem_io_out_0[27:25]; // @[Interconnect.scala 483:23]
  assign Muxn_11_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_4 = io_itrackE_0; // @[Interconnect.scala 475:63]
endmodule
module GIB_11(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire  ConfigMem_clock; // @[Interconnect.scala 463:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 463:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 463:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 463:21]
  wire [27:0] ConfigMem_io_out_0; // @[Interconnect.scala 463:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_6_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_7_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_10_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_11_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_out; // @[Interconnect.scala 473:25]
  wire  _T_1 = 10'h27 == io_cfg_addr[11:2]; // @[Interconnect.scala 464:50]
  reg [31:0] _T_12; // @[Interconnect.scala 477:55]
  reg [31:0] _T_14; // @[Interconnect.scala 477:55]
  reg [31:0] _T_16; // @[Interconnect.scala 477:55]
  reg [31:0] _T_18; // @[Interconnect.scala 477:55]
  ConfigMem_90 ConfigMem ( // @[Interconnect.scala 463:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_148 Muxn ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_out(Muxn_io_out)
  );
  Muxn_148 Muxn_1 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_out(Muxn_1_io_out)
  );
  Muxn_148 Muxn_2 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_in_3(Muxn_2_io_in_3),
    .io_out(Muxn_2_io_out)
  );
  Muxn_148 Muxn_3 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_in_3(Muxn_3_io_in_3),
    .io_out(Muxn_3_io_out)
  );
  Muxn_148 Muxn_4 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_in_3(Muxn_4_io_in_3),
    .io_out(Muxn_4_io_out)
  );
  Muxn_148 Muxn_5 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_in_3(Muxn_5_io_in_3),
    .io_out(Muxn_5_io_out)
  );
  Muxn_148 Muxn_6 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_out(Muxn_6_io_out)
  );
  Muxn_148 Muxn_7 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_out(Muxn_7_io_out)
  );
  Muxn_147 Muxn_8 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_147 Muxn_9 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  Muxn_147 Muxn_10 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_10_io_config),
    .io_in_0(Muxn_10_io_in_0),
    .io_in_1(Muxn_10_io_in_1),
    .io_in_2(Muxn_10_io_in_2),
    .io_in_3(Muxn_10_io_in_3),
    .io_in_4(Muxn_10_io_in_4),
    .io_out(Muxn_10_io_out)
  );
  Muxn_147 Muxn_11 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_11_io_config),
    .io_in_0(Muxn_11_io_in_0),
    .io_in_1(Muxn_11_io_in_1),
    .io_in_2(Muxn_11_io_in_2),
    .io_in_3(Muxn_11_io_in_3),
    .io_in_4(Muxn_11_io_in_4),
    .io_out(Muxn_11_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNE_0 = Muxn_2_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinNE_1 = Muxn_3_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinSE_0 = Muxn_4_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSE_1 = Muxn_5_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSW_0 = Muxn_6_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_ipinSW_1 = Muxn_7_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_otrackW_0 = _T_12; // @[Interconnect.scala 430:21 Interconnect.scala 477:45]
  assign io_otrackN_0 = _T_14; // @[Interconnect.scala 431:21 Interconnect.scala 477:45]
  assign io_otrackE_0 = _T_16; // @[Interconnect.scala 432:21 Interconnect.scala 477:45]
  assign io_otrackS_0 = _T_18; // @[Interconnect.scala 433:21 Interconnect.scala 477:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 464:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 466:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 483:23]
  assign Muxn_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 483:23]
  assign Muxn_1_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 483:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 483:23]
  assign Muxn_3_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 483:23]
  assign Muxn_4_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 483:23]
  assign Muxn_5_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[13:12]; // @[Interconnect.scala 483:23]
  assign Muxn_6_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[15:14]; // @[Interconnect.scala 483:23]
  assign Muxn_7_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[18:16]; // @[Interconnect.scala 483:23]
  assign Muxn_8_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[21:19]; // @[Interconnect.scala 483:23]
  assign Muxn_9_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_config = ConfigMem_io_out_0[24:22]; // @[Interconnect.scala 483:23]
  assign Muxn_10_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_config = ConfigMem_io_out_0[27:25]; // @[Interconnect.scala 483:23]
  assign Muxn_11_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_4 = io_itrackE_0; // @[Interconnect.scala 475:63]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_12 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  _T_14 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  _T_16 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  _T_18 = _RAND_3[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_12 <= Muxn_8_io_out;
    _T_14 <= Muxn_9_io_out;
    _T_16 <= Muxn_10_io_out;
    _T_18 <= Muxn_11_io_out;
  end
endmodule
module GIB_12(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
  wire  ConfigMem_clock; // @[Interconnect.scala 463:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 463:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 463:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 463:21]
  wire [27:0] ConfigMem_io_out_0; // @[Interconnect.scala 463:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_6_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_7_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_10_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_11_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_out; // @[Interconnect.scala 473:25]
  wire  _T_1 = 10'h28 == io_cfg_addr[11:2]; // @[Interconnect.scala 464:50]
  ConfigMem_90 ConfigMem ( // @[Interconnect.scala 463:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_148 Muxn ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_out(Muxn_io_out)
  );
  Muxn_148 Muxn_1 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_out(Muxn_1_io_out)
  );
  Muxn_148 Muxn_2 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_in_3(Muxn_2_io_in_3),
    .io_out(Muxn_2_io_out)
  );
  Muxn_148 Muxn_3 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_in_3(Muxn_3_io_in_3),
    .io_out(Muxn_3_io_out)
  );
  Muxn_148 Muxn_4 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_in_3(Muxn_4_io_in_3),
    .io_out(Muxn_4_io_out)
  );
  Muxn_148 Muxn_5 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_in_3(Muxn_5_io_in_3),
    .io_out(Muxn_5_io_out)
  );
  Muxn_148 Muxn_6 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_out(Muxn_6_io_out)
  );
  Muxn_148 Muxn_7 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_out(Muxn_7_io_out)
  );
  Muxn_147 Muxn_8 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_147 Muxn_9 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  Muxn_147 Muxn_10 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_10_io_config),
    .io_in_0(Muxn_10_io_in_0),
    .io_in_1(Muxn_10_io_in_1),
    .io_in_2(Muxn_10_io_in_2),
    .io_in_3(Muxn_10_io_in_3),
    .io_in_4(Muxn_10_io_in_4),
    .io_out(Muxn_10_io_out)
  );
  Muxn_147 Muxn_11 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_11_io_config),
    .io_in_0(Muxn_11_io_in_0),
    .io_in_1(Muxn_11_io_in_1),
    .io_in_2(Muxn_11_io_in_2),
    .io_in_3(Muxn_11_io_in_3),
    .io_in_4(Muxn_11_io_in_4),
    .io_out(Muxn_11_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNE_0 = Muxn_2_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinNE_1 = Muxn_3_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinSE_0 = Muxn_4_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSE_1 = Muxn_5_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSW_0 = Muxn_6_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_ipinSW_1 = Muxn_7_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_otrackW_0 = Muxn_8_io_out; // @[Interconnect.scala 430:21 Interconnect.scala 479:45]
  assign io_otrackN_0 = Muxn_9_io_out; // @[Interconnect.scala 431:21 Interconnect.scala 479:45]
  assign io_otrackE_0 = Muxn_10_io_out; // @[Interconnect.scala 432:21 Interconnect.scala 479:45]
  assign io_otrackS_0 = Muxn_11_io_out; // @[Interconnect.scala 433:21 Interconnect.scala 479:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 464:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 466:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 483:23]
  assign Muxn_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 483:23]
  assign Muxn_1_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 483:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 483:23]
  assign Muxn_3_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 483:23]
  assign Muxn_4_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 483:23]
  assign Muxn_5_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[13:12]; // @[Interconnect.scala 483:23]
  assign Muxn_6_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[15:14]; // @[Interconnect.scala 483:23]
  assign Muxn_7_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[18:16]; // @[Interconnect.scala 483:23]
  assign Muxn_8_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[21:19]; // @[Interconnect.scala 483:23]
  assign Muxn_9_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_config = ConfigMem_io_out_0[24:22]; // @[Interconnect.scala 483:23]
  assign Muxn_10_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_config = ConfigMem_io_out_0[27:25]; // @[Interconnect.scala 483:23]
  assign Muxn_11_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_4 = io_itrackE_0; // @[Interconnect.scala 475:63]
endmodule
module GIB_13(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire  ConfigMem_clock; // @[Interconnect.scala 463:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 463:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 463:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 463:21]
  wire [27:0] ConfigMem_io_out_0; // @[Interconnect.scala 463:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_6_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_7_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_10_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_11_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_out; // @[Interconnect.scala 473:25]
  wire  _T_1 = 10'h29 == io_cfg_addr[11:2]; // @[Interconnect.scala 464:50]
  reg [31:0] _T_12; // @[Interconnect.scala 477:55]
  reg [31:0] _T_14; // @[Interconnect.scala 477:55]
  reg [31:0] _T_16; // @[Interconnect.scala 477:55]
  reg [31:0] _T_18; // @[Interconnect.scala 477:55]
  ConfigMem_90 ConfigMem ( // @[Interconnect.scala 463:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_148 Muxn ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_out(Muxn_io_out)
  );
  Muxn_148 Muxn_1 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_out(Muxn_1_io_out)
  );
  Muxn_148 Muxn_2 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_in_3(Muxn_2_io_in_3),
    .io_out(Muxn_2_io_out)
  );
  Muxn_148 Muxn_3 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_in_3(Muxn_3_io_in_3),
    .io_out(Muxn_3_io_out)
  );
  Muxn_148 Muxn_4 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_in_3(Muxn_4_io_in_3),
    .io_out(Muxn_4_io_out)
  );
  Muxn_148 Muxn_5 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_in_3(Muxn_5_io_in_3),
    .io_out(Muxn_5_io_out)
  );
  Muxn_148 Muxn_6 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_out(Muxn_6_io_out)
  );
  Muxn_148 Muxn_7 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_out(Muxn_7_io_out)
  );
  Muxn_147 Muxn_8 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_147 Muxn_9 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  Muxn_147 Muxn_10 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_10_io_config),
    .io_in_0(Muxn_10_io_in_0),
    .io_in_1(Muxn_10_io_in_1),
    .io_in_2(Muxn_10_io_in_2),
    .io_in_3(Muxn_10_io_in_3),
    .io_in_4(Muxn_10_io_in_4),
    .io_out(Muxn_10_io_out)
  );
  Muxn_147 Muxn_11 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_11_io_config),
    .io_in_0(Muxn_11_io_in_0),
    .io_in_1(Muxn_11_io_in_1),
    .io_in_2(Muxn_11_io_in_2),
    .io_in_3(Muxn_11_io_in_3),
    .io_in_4(Muxn_11_io_in_4),
    .io_out(Muxn_11_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNE_0 = Muxn_2_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinNE_1 = Muxn_3_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinSE_0 = Muxn_4_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSE_1 = Muxn_5_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSW_0 = Muxn_6_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_ipinSW_1 = Muxn_7_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_otrackW_0 = _T_12; // @[Interconnect.scala 430:21 Interconnect.scala 477:45]
  assign io_otrackN_0 = _T_14; // @[Interconnect.scala 431:21 Interconnect.scala 477:45]
  assign io_otrackE_0 = _T_16; // @[Interconnect.scala 432:21 Interconnect.scala 477:45]
  assign io_otrackS_0 = _T_18; // @[Interconnect.scala 433:21 Interconnect.scala 477:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 464:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 466:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 483:23]
  assign Muxn_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 483:23]
  assign Muxn_1_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 483:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 483:23]
  assign Muxn_3_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 483:23]
  assign Muxn_4_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 483:23]
  assign Muxn_5_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[13:12]; // @[Interconnect.scala 483:23]
  assign Muxn_6_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[15:14]; // @[Interconnect.scala 483:23]
  assign Muxn_7_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[18:16]; // @[Interconnect.scala 483:23]
  assign Muxn_8_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[21:19]; // @[Interconnect.scala 483:23]
  assign Muxn_9_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_config = ConfigMem_io_out_0[24:22]; // @[Interconnect.scala 483:23]
  assign Muxn_10_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_config = ConfigMem_io_out_0[27:25]; // @[Interconnect.scala 483:23]
  assign Muxn_11_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_4 = io_itrackE_0; // @[Interconnect.scala 475:63]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_12 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  _T_14 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  _T_16 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  _T_18 = _RAND_3[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_12 <= Muxn_8_io_out;
    _T_14 <= Muxn_9_io_out;
    _T_16 <= Muxn_10_io_out;
    _T_18 <= Muxn_11_io_out;
  end
endmodule
module GIB_14(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
  wire  ConfigMem_clock; // @[Interconnect.scala 463:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 463:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 463:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 463:21]
  wire [27:0] ConfigMem_io_out_0; // @[Interconnect.scala 463:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_6_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_7_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_10_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_11_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_out; // @[Interconnect.scala 473:25]
  wire  _T_1 = 10'h2a == io_cfg_addr[11:2]; // @[Interconnect.scala 464:50]
  ConfigMem_90 ConfigMem ( // @[Interconnect.scala 463:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_148 Muxn ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_out(Muxn_io_out)
  );
  Muxn_148 Muxn_1 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_out(Muxn_1_io_out)
  );
  Muxn_148 Muxn_2 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_in_3(Muxn_2_io_in_3),
    .io_out(Muxn_2_io_out)
  );
  Muxn_148 Muxn_3 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_in_3(Muxn_3_io_in_3),
    .io_out(Muxn_3_io_out)
  );
  Muxn_148 Muxn_4 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_in_3(Muxn_4_io_in_3),
    .io_out(Muxn_4_io_out)
  );
  Muxn_148 Muxn_5 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_in_3(Muxn_5_io_in_3),
    .io_out(Muxn_5_io_out)
  );
  Muxn_148 Muxn_6 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_out(Muxn_6_io_out)
  );
  Muxn_148 Muxn_7 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_out(Muxn_7_io_out)
  );
  Muxn_147 Muxn_8 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_147 Muxn_9 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  Muxn_147 Muxn_10 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_10_io_config),
    .io_in_0(Muxn_10_io_in_0),
    .io_in_1(Muxn_10_io_in_1),
    .io_in_2(Muxn_10_io_in_2),
    .io_in_3(Muxn_10_io_in_3),
    .io_in_4(Muxn_10_io_in_4),
    .io_out(Muxn_10_io_out)
  );
  Muxn_147 Muxn_11 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_11_io_config),
    .io_in_0(Muxn_11_io_in_0),
    .io_in_1(Muxn_11_io_in_1),
    .io_in_2(Muxn_11_io_in_2),
    .io_in_3(Muxn_11_io_in_3),
    .io_in_4(Muxn_11_io_in_4),
    .io_out(Muxn_11_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNE_0 = Muxn_2_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinNE_1 = Muxn_3_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinSE_0 = Muxn_4_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSE_1 = Muxn_5_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSW_0 = Muxn_6_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_ipinSW_1 = Muxn_7_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_otrackW_0 = Muxn_8_io_out; // @[Interconnect.scala 430:21 Interconnect.scala 479:45]
  assign io_otrackN_0 = Muxn_9_io_out; // @[Interconnect.scala 431:21 Interconnect.scala 479:45]
  assign io_otrackE_0 = Muxn_10_io_out; // @[Interconnect.scala 432:21 Interconnect.scala 479:45]
  assign io_otrackS_0 = Muxn_11_io_out; // @[Interconnect.scala 433:21 Interconnect.scala 479:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 464:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 466:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 483:23]
  assign Muxn_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 483:23]
  assign Muxn_1_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 483:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 483:23]
  assign Muxn_3_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 483:23]
  assign Muxn_4_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 483:23]
  assign Muxn_5_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[13:12]; // @[Interconnect.scala 483:23]
  assign Muxn_6_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[15:14]; // @[Interconnect.scala 483:23]
  assign Muxn_7_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[18:16]; // @[Interconnect.scala 483:23]
  assign Muxn_8_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[21:19]; // @[Interconnect.scala 483:23]
  assign Muxn_9_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_config = ConfigMem_io_out_0[24:22]; // @[Interconnect.scala 483:23]
  assign Muxn_10_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_config = ConfigMem_io_out_0[27:25]; // @[Interconnect.scala 483:23]
  assign Muxn_11_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_4 = io_itrackE_0; // @[Interconnect.scala 475:63]
endmodule
module GIB_15(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire  ConfigMem_clock; // @[Interconnect.scala 463:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 463:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 463:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 463:21]
  wire [27:0] ConfigMem_io_out_0; // @[Interconnect.scala 463:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_6_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_7_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_10_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_11_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_out; // @[Interconnect.scala 473:25]
  wire  _T_1 = 10'h2b == io_cfg_addr[11:2]; // @[Interconnect.scala 464:50]
  reg [31:0] _T_12; // @[Interconnect.scala 477:55]
  reg [31:0] _T_14; // @[Interconnect.scala 477:55]
  reg [31:0] _T_16; // @[Interconnect.scala 477:55]
  reg [31:0] _T_18; // @[Interconnect.scala 477:55]
  ConfigMem_90 ConfigMem ( // @[Interconnect.scala 463:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_148 Muxn ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_out(Muxn_io_out)
  );
  Muxn_148 Muxn_1 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_out(Muxn_1_io_out)
  );
  Muxn_148 Muxn_2 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_in_3(Muxn_2_io_in_3),
    .io_out(Muxn_2_io_out)
  );
  Muxn_148 Muxn_3 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_in_3(Muxn_3_io_in_3),
    .io_out(Muxn_3_io_out)
  );
  Muxn_148 Muxn_4 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_in_3(Muxn_4_io_in_3),
    .io_out(Muxn_4_io_out)
  );
  Muxn_148 Muxn_5 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_in_3(Muxn_5_io_in_3),
    .io_out(Muxn_5_io_out)
  );
  Muxn_148 Muxn_6 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_out(Muxn_6_io_out)
  );
  Muxn_148 Muxn_7 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_out(Muxn_7_io_out)
  );
  Muxn_147 Muxn_8 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_147 Muxn_9 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  Muxn_147 Muxn_10 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_10_io_config),
    .io_in_0(Muxn_10_io_in_0),
    .io_in_1(Muxn_10_io_in_1),
    .io_in_2(Muxn_10_io_in_2),
    .io_in_3(Muxn_10_io_in_3),
    .io_in_4(Muxn_10_io_in_4),
    .io_out(Muxn_10_io_out)
  );
  Muxn_147 Muxn_11 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_11_io_config),
    .io_in_0(Muxn_11_io_in_0),
    .io_in_1(Muxn_11_io_in_1),
    .io_in_2(Muxn_11_io_in_2),
    .io_in_3(Muxn_11_io_in_3),
    .io_in_4(Muxn_11_io_in_4),
    .io_out(Muxn_11_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNE_0 = Muxn_2_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinNE_1 = Muxn_3_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinSE_0 = Muxn_4_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSE_1 = Muxn_5_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSW_0 = Muxn_6_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_ipinSW_1 = Muxn_7_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_otrackW_0 = _T_12; // @[Interconnect.scala 430:21 Interconnect.scala 477:45]
  assign io_otrackN_0 = _T_14; // @[Interconnect.scala 431:21 Interconnect.scala 477:45]
  assign io_otrackE_0 = _T_16; // @[Interconnect.scala 432:21 Interconnect.scala 477:45]
  assign io_otrackS_0 = _T_18; // @[Interconnect.scala 433:21 Interconnect.scala 477:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 464:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 466:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 483:23]
  assign Muxn_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 483:23]
  assign Muxn_1_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 483:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 483:23]
  assign Muxn_3_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 483:23]
  assign Muxn_4_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 483:23]
  assign Muxn_5_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[13:12]; // @[Interconnect.scala 483:23]
  assign Muxn_6_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[15:14]; // @[Interconnect.scala 483:23]
  assign Muxn_7_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[18:16]; // @[Interconnect.scala 483:23]
  assign Muxn_8_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[21:19]; // @[Interconnect.scala 483:23]
  assign Muxn_9_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_config = ConfigMem_io_out_0[24:22]; // @[Interconnect.scala 483:23]
  assign Muxn_10_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_config = ConfigMem_io_out_0[27:25]; // @[Interconnect.scala 483:23]
  assign Muxn_11_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_4 = io_itrackE_0; // @[Interconnect.scala 475:63]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_12 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  _T_14 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  _T_16 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  _T_18 = _RAND_3[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_12 <= Muxn_8_io_out;
    _T_14 <= Muxn_9_io_out;
    _T_16 <= Muxn_10_io_out;
    _T_18 <= Muxn_11_io_out;
  end
endmodule
module GIB_16(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
  wire  ConfigMem_clock; // @[Interconnect.scala 463:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 463:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 463:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 463:21]
  wire [27:0] ConfigMem_io_out_0; // @[Interconnect.scala 463:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_6_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_7_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_10_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_11_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_out; // @[Interconnect.scala 473:25]
  wire  _T_1 = 10'h2c == io_cfg_addr[11:2]; // @[Interconnect.scala 464:50]
  ConfigMem_90 ConfigMem ( // @[Interconnect.scala 463:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_148 Muxn ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_out(Muxn_io_out)
  );
  Muxn_148 Muxn_1 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_out(Muxn_1_io_out)
  );
  Muxn_148 Muxn_2 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_in_3(Muxn_2_io_in_3),
    .io_out(Muxn_2_io_out)
  );
  Muxn_148 Muxn_3 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_in_3(Muxn_3_io_in_3),
    .io_out(Muxn_3_io_out)
  );
  Muxn_148 Muxn_4 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_in_3(Muxn_4_io_in_3),
    .io_out(Muxn_4_io_out)
  );
  Muxn_148 Muxn_5 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_in_3(Muxn_5_io_in_3),
    .io_out(Muxn_5_io_out)
  );
  Muxn_148 Muxn_6 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_out(Muxn_6_io_out)
  );
  Muxn_148 Muxn_7 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_out(Muxn_7_io_out)
  );
  Muxn_147 Muxn_8 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_147 Muxn_9 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  Muxn_147 Muxn_10 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_10_io_config),
    .io_in_0(Muxn_10_io_in_0),
    .io_in_1(Muxn_10_io_in_1),
    .io_in_2(Muxn_10_io_in_2),
    .io_in_3(Muxn_10_io_in_3),
    .io_in_4(Muxn_10_io_in_4),
    .io_out(Muxn_10_io_out)
  );
  Muxn_147 Muxn_11 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_11_io_config),
    .io_in_0(Muxn_11_io_in_0),
    .io_in_1(Muxn_11_io_in_1),
    .io_in_2(Muxn_11_io_in_2),
    .io_in_3(Muxn_11_io_in_3),
    .io_in_4(Muxn_11_io_in_4),
    .io_out(Muxn_11_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNE_0 = Muxn_2_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinNE_1 = Muxn_3_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinSE_0 = Muxn_4_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSE_1 = Muxn_5_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSW_0 = Muxn_6_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_ipinSW_1 = Muxn_7_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_otrackW_0 = Muxn_8_io_out; // @[Interconnect.scala 430:21 Interconnect.scala 479:45]
  assign io_otrackN_0 = Muxn_9_io_out; // @[Interconnect.scala 431:21 Interconnect.scala 479:45]
  assign io_otrackE_0 = Muxn_10_io_out; // @[Interconnect.scala 432:21 Interconnect.scala 479:45]
  assign io_otrackS_0 = Muxn_11_io_out; // @[Interconnect.scala 433:21 Interconnect.scala 479:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 464:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 466:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 483:23]
  assign Muxn_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 483:23]
  assign Muxn_1_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 483:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 483:23]
  assign Muxn_3_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 483:23]
  assign Muxn_4_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 483:23]
  assign Muxn_5_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[13:12]; // @[Interconnect.scala 483:23]
  assign Muxn_6_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[15:14]; // @[Interconnect.scala 483:23]
  assign Muxn_7_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[18:16]; // @[Interconnect.scala 483:23]
  assign Muxn_8_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[21:19]; // @[Interconnect.scala 483:23]
  assign Muxn_9_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_config = ConfigMem_io_out_0[24:22]; // @[Interconnect.scala 483:23]
  assign Muxn_10_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_config = ConfigMem_io_out_0[27:25]; // @[Interconnect.scala 483:23]
  assign Muxn_11_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_4 = io_itrackE_0; // @[Interconnect.scala 475:63]
endmodule
module GIB_17(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire  ConfigMem_clock; // @[Interconnect.scala 463:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 463:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 463:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 463:21]
  wire [14:0] ConfigMem_io_out_0; // @[Interconnect.scala 463:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 473:25]
  wire  Muxn_2_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 473:25]
  wire  Muxn_3_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_6_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_7_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 473:25]
  wire  _T_1 = 10'h2d == io_cfg_addr[11:2]; // @[Interconnect.scala 464:50]
  reg [31:0] _T_8; // @[Interconnect.scala 477:55]
  reg [31:0] _T_10; // @[Interconnect.scala 477:55]
  reg [31:0] _T_14; // @[Interconnect.scala 477:55]
  ConfigMem_89 ConfigMem ( // @[Interconnect.scala 463:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_145 Muxn ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_out(Muxn_io_out)
  );
  Muxn_145 Muxn_1 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_out(Muxn_1_io_out)
  );
  Muxn Muxn_2 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_out(Muxn_2_io_out)
  );
  Muxn Muxn_3 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_out(Muxn_3_io_out)
  );
  Muxn_145 Muxn_4 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_out(Muxn_4_io_out)
  );
  Muxn_148 Muxn_5 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_in_3(Muxn_5_io_in_3),
    .io_out(Muxn_5_io_out)
  );
  Muxn_147 Muxn_6 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_in_4(Muxn_6_io_in_4),
    .io_out(Muxn_6_io_out)
  );
  Muxn_148 Muxn_7 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_out(Muxn_7_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinSW_0 = Muxn_2_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_ipinSW_1 = Muxn_3_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_otrackW_0 = _T_8; // @[Interconnect.scala 430:21 Interconnect.scala 477:45]
  assign io_otrackN_0 = _T_10; // @[Interconnect.scala 431:21 Interconnect.scala 477:45]
  assign io_otrackS_0 = _T_14; // @[Interconnect.scala 433:21 Interconnect.scala 477:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 464:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 466:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 483:23]
  assign Muxn_io_in_0 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_1 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_2 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 483:23]
  assign Muxn_1_io_in_0 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_1 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_2 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[4]; // @[Interconnect.scala 483:23]
  assign Muxn_2_io_in_0 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_1 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[5]; // @[Interconnect.scala 483:23]
  assign Muxn_3_io_in_0 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_1 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 483:23]
  assign Muxn_4_io_in_0 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_1 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_2 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 483:23]
  assign Muxn_5_io_in_0 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_1 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_2 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[12:10]; // @[Interconnect.scala 483:23]
  assign Muxn_6_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[14:13]; // @[Interconnect.scala 483:23]
  assign Muxn_7_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_1 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_3 = 32'h0; // @[Interconnect.scala 475:63]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_8 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  _T_10 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  _T_14 = _RAND_2[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_8 <= Muxn_4_io_out;
    _T_10 <= Muxn_5_io_out;
    _T_14 <= Muxn_7_io_out;
  end
endmodule
module GIB_18(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
  wire  ConfigMem_clock; // @[Interconnect.scala 463:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 463:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 463:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 463:21]
  wire [14:0] ConfigMem_io_out_0; // @[Interconnect.scala 463:21]
  wire  Muxn_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 473:25]
  wire  Muxn_1_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_4_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_6_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_7_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 473:25]
  wire  _T_1 = 10'h37 == io_cfg_addr[11:2]; // @[Interconnect.scala 464:50]
  ConfigMem_89 ConfigMem ( // @[Interconnect.scala 463:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn Muxn ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_out(Muxn_io_out)
  );
  Muxn Muxn_1 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_out(Muxn_1_io_out)
  );
  Muxn_145 Muxn_2 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_out(Muxn_2_io_out)
  );
  Muxn_145 Muxn_3 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_out(Muxn_3_io_out)
  );
  Muxn_147 Muxn_4 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_in_3(Muxn_4_io_in_3),
    .io_in_4(Muxn_4_io_in_4),
    .io_out(Muxn_4_io_out)
  );
  Muxn_148 Muxn_5 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_in_3(Muxn_5_io_in_3),
    .io_out(Muxn_5_io_out)
  );
  Muxn_145 Muxn_6 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_out(Muxn_6_io_out)
  );
  Muxn_148 Muxn_7 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_out(Muxn_7_io_out)
  );
  assign io_ipinNE_0 = Muxn_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinNE_1 = Muxn_1_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinSE_0 = Muxn_2_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSE_1 = Muxn_3_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_otrackN_0 = Muxn_5_io_out; // @[Interconnect.scala 431:21 Interconnect.scala 479:45]
  assign io_otrackE_0 = Muxn_6_io_out; // @[Interconnect.scala 432:21 Interconnect.scala 479:45]
  assign io_otrackS_0 = Muxn_7_io_out; // @[Interconnect.scala 433:21 Interconnect.scala 479:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 464:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 466:21]
  assign Muxn_io_config = ConfigMem_io_out_0[0]; // @[Interconnect.scala 483:23]
  assign Muxn_io_in_0 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_1 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[1]; // @[Interconnect.scala 483:23]
  assign Muxn_1_io_in_0 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_1 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 483:23]
  assign Muxn_2_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_1 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 483:23]
  assign Muxn_3_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_1 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[8:6]; // @[Interconnect.scala 483:23]
  assign Muxn_4_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[10:9]; // @[Interconnect.scala 483:23]
  assign Muxn_5_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_1 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[12:11]; // @[Interconnect.scala 483:23]
  assign Muxn_6_io_in_0 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_1 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_2 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[14:13]; // @[Interconnect.scala 483:23]
  assign Muxn_7_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_1 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
endmodule
module GIB_19(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire  ConfigMem_clock; // @[Interconnect.scala 463:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 463:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 463:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 463:21]
  wire [27:0] ConfigMem_io_out_0; // @[Interconnect.scala 463:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_6_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_7_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_10_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_11_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_out; // @[Interconnect.scala 473:25]
  wire  _T_1 = 10'h38 == io_cfg_addr[11:2]; // @[Interconnect.scala 464:50]
  reg [31:0] _T_12; // @[Interconnect.scala 477:55]
  reg [31:0] _T_14; // @[Interconnect.scala 477:55]
  reg [31:0] _T_16; // @[Interconnect.scala 477:55]
  reg [31:0] _T_18; // @[Interconnect.scala 477:55]
  ConfigMem_90 ConfigMem ( // @[Interconnect.scala 463:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_148 Muxn ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_out(Muxn_io_out)
  );
  Muxn_148 Muxn_1 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_out(Muxn_1_io_out)
  );
  Muxn_148 Muxn_2 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_in_3(Muxn_2_io_in_3),
    .io_out(Muxn_2_io_out)
  );
  Muxn_148 Muxn_3 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_in_3(Muxn_3_io_in_3),
    .io_out(Muxn_3_io_out)
  );
  Muxn_148 Muxn_4 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_in_3(Muxn_4_io_in_3),
    .io_out(Muxn_4_io_out)
  );
  Muxn_148 Muxn_5 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_in_3(Muxn_5_io_in_3),
    .io_out(Muxn_5_io_out)
  );
  Muxn_148 Muxn_6 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_out(Muxn_6_io_out)
  );
  Muxn_148 Muxn_7 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_out(Muxn_7_io_out)
  );
  Muxn_147 Muxn_8 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_147 Muxn_9 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  Muxn_147 Muxn_10 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_10_io_config),
    .io_in_0(Muxn_10_io_in_0),
    .io_in_1(Muxn_10_io_in_1),
    .io_in_2(Muxn_10_io_in_2),
    .io_in_3(Muxn_10_io_in_3),
    .io_in_4(Muxn_10_io_in_4),
    .io_out(Muxn_10_io_out)
  );
  Muxn_147 Muxn_11 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_11_io_config),
    .io_in_0(Muxn_11_io_in_0),
    .io_in_1(Muxn_11_io_in_1),
    .io_in_2(Muxn_11_io_in_2),
    .io_in_3(Muxn_11_io_in_3),
    .io_in_4(Muxn_11_io_in_4),
    .io_out(Muxn_11_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNE_0 = Muxn_2_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinNE_1 = Muxn_3_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinSE_0 = Muxn_4_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSE_1 = Muxn_5_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSW_0 = Muxn_6_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_ipinSW_1 = Muxn_7_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_otrackW_0 = _T_12; // @[Interconnect.scala 430:21 Interconnect.scala 477:45]
  assign io_otrackN_0 = _T_14; // @[Interconnect.scala 431:21 Interconnect.scala 477:45]
  assign io_otrackE_0 = _T_16; // @[Interconnect.scala 432:21 Interconnect.scala 477:45]
  assign io_otrackS_0 = _T_18; // @[Interconnect.scala 433:21 Interconnect.scala 477:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 464:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 466:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 483:23]
  assign Muxn_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 483:23]
  assign Muxn_1_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 483:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 483:23]
  assign Muxn_3_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 483:23]
  assign Muxn_4_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 483:23]
  assign Muxn_5_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[13:12]; // @[Interconnect.scala 483:23]
  assign Muxn_6_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[15:14]; // @[Interconnect.scala 483:23]
  assign Muxn_7_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[18:16]; // @[Interconnect.scala 483:23]
  assign Muxn_8_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[21:19]; // @[Interconnect.scala 483:23]
  assign Muxn_9_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_config = ConfigMem_io_out_0[24:22]; // @[Interconnect.scala 483:23]
  assign Muxn_10_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_config = ConfigMem_io_out_0[27:25]; // @[Interconnect.scala 483:23]
  assign Muxn_11_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_4 = io_itrackE_0; // @[Interconnect.scala 475:63]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_12 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  _T_14 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  _T_16 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  _T_18 = _RAND_3[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_12 <= Muxn_8_io_out;
    _T_14 <= Muxn_9_io_out;
    _T_16 <= Muxn_10_io_out;
    _T_18 <= Muxn_11_io_out;
  end
endmodule
module GIB_20(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
  wire  ConfigMem_clock; // @[Interconnect.scala 463:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 463:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 463:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 463:21]
  wire [27:0] ConfigMem_io_out_0; // @[Interconnect.scala 463:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_6_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_7_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_10_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_11_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_out; // @[Interconnect.scala 473:25]
  wire  _T_1 = 10'h39 == io_cfg_addr[11:2]; // @[Interconnect.scala 464:50]
  ConfigMem_90 ConfigMem ( // @[Interconnect.scala 463:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_148 Muxn ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_out(Muxn_io_out)
  );
  Muxn_148 Muxn_1 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_out(Muxn_1_io_out)
  );
  Muxn_148 Muxn_2 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_in_3(Muxn_2_io_in_3),
    .io_out(Muxn_2_io_out)
  );
  Muxn_148 Muxn_3 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_in_3(Muxn_3_io_in_3),
    .io_out(Muxn_3_io_out)
  );
  Muxn_148 Muxn_4 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_in_3(Muxn_4_io_in_3),
    .io_out(Muxn_4_io_out)
  );
  Muxn_148 Muxn_5 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_in_3(Muxn_5_io_in_3),
    .io_out(Muxn_5_io_out)
  );
  Muxn_148 Muxn_6 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_out(Muxn_6_io_out)
  );
  Muxn_148 Muxn_7 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_out(Muxn_7_io_out)
  );
  Muxn_147 Muxn_8 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_147 Muxn_9 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  Muxn_147 Muxn_10 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_10_io_config),
    .io_in_0(Muxn_10_io_in_0),
    .io_in_1(Muxn_10_io_in_1),
    .io_in_2(Muxn_10_io_in_2),
    .io_in_3(Muxn_10_io_in_3),
    .io_in_4(Muxn_10_io_in_4),
    .io_out(Muxn_10_io_out)
  );
  Muxn_147 Muxn_11 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_11_io_config),
    .io_in_0(Muxn_11_io_in_0),
    .io_in_1(Muxn_11_io_in_1),
    .io_in_2(Muxn_11_io_in_2),
    .io_in_3(Muxn_11_io_in_3),
    .io_in_4(Muxn_11_io_in_4),
    .io_out(Muxn_11_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNE_0 = Muxn_2_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinNE_1 = Muxn_3_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinSE_0 = Muxn_4_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSE_1 = Muxn_5_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSW_0 = Muxn_6_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_ipinSW_1 = Muxn_7_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_otrackW_0 = Muxn_8_io_out; // @[Interconnect.scala 430:21 Interconnect.scala 479:45]
  assign io_otrackN_0 = Muxn_9_io_out; // @[Interconnect.scala 431:21 Interconnect.scala 479:45]
  assign io_otrackE_0 = Muxn_10_io_out; // @[Interconnect.scala 432:21 Interconnect.scala 479:45]
  assign io_otrackS_0 = Muxn_11_io_out; // @[Interconnect.scala 433:21 Interconnect.scala 479:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 464:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 466:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 483:23]
  assign Muxn_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 483:23]
  assign Muxn_1_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 483:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 483:23]
  assign Muxn_3_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 483:23]
  assign Muxn_4_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 483:23]
  assign Muxn_5_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[13:12]; // @[Interconnect.scala 483:23]
  assign Muxn_6_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[15:14]; // @[Interconnect.scala 483:23]
  assign Muxn_7_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[18:16]; // @[Interconnect.scala 483:23]
  assign Muxn_8_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[21:19]; // @[Interconnect.scala 483:23]
  assign Muxn_9_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_config = ConfigMem_io_out_0[24:22]; // @[Interconnect.scala 483:23]
  assign Muxn_10_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_config = ConfigMem_io_out_0[27:25]; // @[Interconnect.scala 483:23]
  assign Muxn_11_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_4 = io_itrackE_0; // @[Interconnect.scala 475:63]
endmodule
module GIB_21(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire  ConfigMem_clock; // @[Interconnect.scala 463:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 463:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 463:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 463:21]
  wire [27:0] ConfigMem_io_out_0; // @[Interconnect.scala 463:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_6_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_7_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_10_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_11_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_out; // @[Interconnect.scala 473:25]
  wire  _T_1 = 10'h3a == io_cfg_addr[11:2]; // @[Interconnect.scala 464:50]
  reg [31:0] _T_12; // @[Interconnect.scala 477:55]
  reg [31:0] _T_14; // @[Interconnect.scala 477:55]
  reg [31:0] _T_16; // @[Interconnect.scala 477:55]
  reg [31:0] _T_18; // @[Interconnect.scala 477:55]
  ConfigMem_90 ConfigMem ( // @[Interconnect.scala 463:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_148 Muxn ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_out(Muxn_io_out)
  );
  Muxn_148 Muxn_1 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_out(Muxn_1_io_out)
  );
  Muxn_148 Muxn_2 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_in_3(Muxn_2_io_in_3),
    .io_out(Muxn_2_io_out)
  );
  Muxn_148 Muxn_3 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_in_3(Muxn_3_io_in_3),
    .io_out(Muxn_3_io_out)
  );
  Muxn_148 Muxn_4 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_in_3(Muxn_4_io_in_3),
    .io_out(Muxn_4_io_out)
  );
  Muxn_148 Muxn_5 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_in_3(Muxn_5_io_in_3),
    .io_out(Muxn_5_io_out)
  );
  Muxn_148 Muxn_6 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_out(Muxn_6_io_out)
  );
  Muxn_148 Muxn_7 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_out(Muxn_7_io_out)
  );
  Muxn_147 Muxn_8 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_147 Muxn_9 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  Muxn_147 Muxn_10 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_10_io_config),
    .io_in_0(Muxn_10_io_in_0),
    .io_in_1(Muxn_10_io_in_1),
    .io_in_2(Muxn_10_io_in_2),
    .io_in_3(Muxn_10_io_in_3),
    .io_in_4(Muxn_10_io_in_4),
    .io_out(Muxn_10_io_out)
  );
  Muxn_147 Muxn_11 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_11_io_config),
    .io_in_0(Muxn_11_io_in_0),
    .io_in_1(Muxn_11_io_in_1),
    .io_in_2(Muxn_11_io_in_2),
    .io_in_3(Muxn_11_io_in_3),
    .io_in_4(Muxn_11_io_in_4),
    .io_out(Muxn_11_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNE_0 = Muxn_2_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinNE_1 = Muxn_3_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinSE_0 = Muxn_4_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSE_1 = Muxn_5_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSW_0 = Muxn_6_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_ipinSW_1 = Muxn_7_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_otrackW_0 = _T_12; // @[Interconnect.scala 430:21 Interconnect.scala 477:45]
  assign io_otrackN_0 = _T_14; // @[Interconnect.scala 431:21 Interconnect.scala 477:45]
  assign io_otrackE_0 = _T_16; // @[Interconnect.scala 432:21 Interconnect.scala 477:45]
  assign io_otrackS_0 = _T_18; // @[Interconnect.scala 433:21 Interconnect.scala 477:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 464:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 466:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 483:23]
  assign Muxn_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 483:23]
  assign Muxn_1_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 483:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 483:23]
  assign Muxn_3_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 483:23]
  assign Muxn_4_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 483:23]
  assign Muxn_5_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[13:12]; // @[Interconnect.scala 483:23]
  assign Muxn_6_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[15:14]; // @[Interconnect.scala 483:23]
  assign Muxn_7_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[18:16]; // @[Interconnect.scala 483:23]
  assign Muxn_8_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[21:19]; // @[Interconnect.scala 483:23]
  assign Muxn_9_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_config = ConfigMem_io_out_0[24:22]; // @[Interconnect.scala 483:23]
  assign Muxn_10_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_config = ConfigMem_io_out_0[27:25]; // @[Interconnect.scala 483:23]
  assign Muxn_11_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_4 = io_itrackE_0; // @[Interconnect.scala 475:63]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_12 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  _T_14 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  _T_16 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  _T_18 = _RAND_3[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_12 <= Muxn_8_io_out;
    _T_14 <= Muxn_9_io_out;
    _T_16 <= Muxn_10_io_out;
    _T_18 <= Muxn_11_io_out;
  end
endmodule
module GIB_22(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
  wire  ConfigMem_clock; // @[Interconnect.scala 463:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 463:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 463:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 463:21]
  wire [27:0] ConfigMem_io_out_0; // @[Interconnect.scala 463:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_6_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_7_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_10_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_11_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_out; // @[Interconnect.scala 473:25]
  wire  _T_1 = 10'h3b == io_cfg_addr[11:2]; // @[Interconnect.scala 464:50]
  ConfigMem_90 ConfigMem ( // @[Interconnect.scala 463:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_148 Muxn ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_out(Muxn_io_out)
  );
  Muxn_148 Muxn_1 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_out(Muxn_1_io_out)
  );
  Muxn_148 Muxn_2 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_in_3(Muxn_2_io_in_3),
    .io_out(Muxn_2_io_out)
  );
  Muxn_148 Muxn_3 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_in_3(Muxn_3_io_in_3),
    .io_out(Muxn_3_io_out)
  );
  Muxn_148 Muxn_4 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_in_3(Muxn_4_io_in_3),
    .io_out(Muxn_4_io_out)
  );
  Muxn_148 Muxn_5 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_in_3(Muxn_5_io_in_3),
    .io_out(Muxn_5_io_out)
  );
  Muxn_148 Muxn_6 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_out(Muxn_6_io_out)
  );
  Muxn_148 Muxn_7 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_out(Muxn_7_io_out)
  );
  Muxn_147 Muxn_8 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_147 Muxn_9 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  Muxn_147 Muxn_10 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_10_io_config),
    .io_in_0(Muxn_10_io_in_0),
    .io_in_1(Muxn_10_io_in_1),
    .io_in_2(Muxn_10_io_in_2),
    .io_in_3(Muxn_10_io_in_3),
    .io_in_4(Muxn_10_io_in_4),
    .io_out(Muxn_10_io_out)
  );
  Muxn_147 Muxn_11 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_11_io_config),
    .io_in_0(Muxn_11_io_in_0),
    .io_in_1(Muxn_11_io_in_1),
    .io_in_2(Muxn_11_io_in_2),
    .io_in_3(Muxn_11_io_in_3),
    .io_in_4(Muxn_11_io_in_4),
    .io_out(Muxn_11_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNE_0 = Muxn_2_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinNE_1 = Muxn_3_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinSE_0 = Muxn_4_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSE_1 = Muxn_5_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSW_0 = Muxn_6_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_ipinSW_1 = Muxn_7_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_otrackW_0 = Muxn_8_io_out; // @[Interconnect.scala 430:21 Interconnect.scala 479:45]
  assign io_otrackN_0 = Muxn_9_io_out; // @[Interconnect.scala 431:21 Interconnect.scala 479:45]
  assign io_otrackE_0 = Muxn_10_io_out; // @[Interconnect.scala 432:21 Interconnect.scala 479:45]
  assign io_otrackS_0 = Muxn_11_io_out; // @[Interconnect.scala 433:21 Interconnect.scala 479:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 464:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 466:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 483:23]
  assign Muxn_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 483:23]
  assign Muxn_1_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 483:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 483:23]
  assign Muxn_3_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 483:23]
  assign Muxn_4_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 483:23]
  assign Muxn_5_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[13:12]; // @[Interconnect.scala 483:23]
  assign Muxn_6_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[15:14]; // @[Interconnect.scala 483:23]
  assign Muxn_7_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[18:16]; // @[Interconnect.scala 483:23]
  assign Muxn_8_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[21:19]; // @[Interconnect.scala 483:23]
  assign Muxn_9_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_config = ConfigMem_io_out_0[24:22]; // @[Interconnect.scala 483:23]
  assign Muxn_10_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_config = ConfigMem_io_out_0[27:25]; // @[Interconnect.scala 483:23]
  assign Muxn_11_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_4 = io_itrackE_0; // @[Interconnect.scala 475:63]
endmodule
module GIB_23(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire  ConfigMem_clock; // @[Interconnect.scala 463:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 463:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 463:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 463:21]
  wire [27:0] ConfigMem_io_out_0; // @[Interconnect.scala 463:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_6_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_7_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_10_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_11_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_out; // @[Interconnect.scala 473:25]
  wire  _T_1 = 10'h3c == io_cfg_addr[11:2]; // @[Interconnect.scala 464:50]
  reg [31:0] _T_12; // @[Interconnect.scala 477:55]
  reg [31:0] _T_14; // @[Interconnect.scala 477:55]
  reg [31:0] _T_16; // @[Interconnect.scala 477:55]
  reg [31:0] _T_18; // @[Interconnect.scala 477:55]
  ConfigMem_90 ConfigMem ( // @[Interconnect.scala 463:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_148 Muxn ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_out(Muxn_io_out)
  );
  Muxn_148 Muxn_1 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_out(Muxn_1_io_out)
  );
  Muxn_148 Muxn_2 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_in_3(Muxn_2_io_in_3),
    .io_out(Muxn_2_io_out)
  );
  Muxn_148 Muxn_3 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_in_3(Muxn_3_io_in_3),
    .io_out(Muxn_3_io_out)
  );
  Muxn_148 Muxn_4 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_in_3(Muxn_4_io_in_3),
    .io_out(Muxn_4_io_out)
  );
  Muxn_148 Muxn_5 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_in_3(Muxn_5_io_in_3),
    .io_out(Muxn_5_io_out)
  );
  Muxn_148 Muxn_6 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_out(Muxn_6_io_out)
  );
  Muxn_148 Muxn_7 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_out(Muxn_7_io_out)
  );
  Muxn_147 Muxn_8 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_147 Muxn_9 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  Muxn_147 Muxn_10 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_10_io_config),
    .io_in_0(Muxn_10_io_in_0),
    .io_in_1(Muxn_10_io_in_1),
    .io_in_2(Muxn_10_io_in_2),
    .io_in_3(Muxn_10_io_in_3),
    .io_in_4(Muxn_10_io_in_4),
    .io_out(Muxn_10_io_out)
  );
  Muxn_147 Muxn_11 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_11_io_config),
    .io_in_0(Muxn_11_io_in_0),
    .io_in_1(Muxn_11_io_in_1),
    .io_in_2(Muxn_11_io_in_2),
    .io_in_3(Muxn_11_io_in_3),
    .io_in_4(Muxn_11_io_in_4),
    .io_out(Muxn_11_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNE_0 = Muxn_2_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinNE_1 = Muxn_3_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinSE_0 = Muxn_4_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSE_1 = Muxn_5_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSW_0 = Muxn_6_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_ipinSW_1 = Muxn_7_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_otrackW_0 = _T_12; // @[Interconnect.scala 430:21 Interconnect.scala 477:45]
  assign io_otrackN_0 = _T_14; // @[Interconnect.scala 431:21 Interconnect.scala 477:45]
  assign io_otrackE_0 = _T_16; // @[Interconnect.scala 432:21 Interconnect.scala 477:45]
  assign io_otrackS_0 = _T_18; // @[Interconnect.scala 433:21 Interconnect.scala 477:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 464:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 466:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 483:23]
  assign Muxn_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 483:23]
  assign Muxn_1_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 483:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 483:23]
  assign Muxn_3_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 483:23]
  assign Muxn_4_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 483:23]
  assign Muxn_5_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[13:12]; // @[Interconnect.scala 483:23]
  assign Muxn_6_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[15:14]; // @[Interconnect.scala 483:23]
  assign Muxn_7_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[18:16]; // @[Interconnect.scala 483:23]
  assign Muxn_8_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[21:19]; // @[Interconnect.scala 483:23]
  assign Muxn_9_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_config = ConfigMem_io_out_0[24:22]; // @[Interconnect.scala 483:23]
  assign Muxn_10_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_config = ConfigMem_io_out_0[27:25]; // @[Interconnect.scala 483:23]
  assign Muxn_11_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_4 = io_itrackE_0; // @[Interconnect.scala 475:63]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_12 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  _T_14 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  _T_16 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  _T_18 = _RAND_3[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_12 <= Muxn_8_io_out;
    _T_14 <= Muxn_9_io_out;
    _T_16 <= Muxn_10_io_out;
    _T_18 <= Muxn_11_io_out;
  end
endmodule
module GIB_24(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
  wire  ConfigMem_clock; // @[Interconnect.scala 463:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 463:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 463:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 463:21]
  wire [27:0] ConfigMem_io_out_0; // @[Interconnect.scala 463:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_6_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_7_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_10_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_11_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_out; // @[Interconnect.scala 473:25]
  wire  _T_1 = 10'h3d == io_cfg_addr[11:2]; // @[Interconnect.scala 464:50]
  ConfigMem_90 ConfigMem ( // @[Interconnect.scala 463:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_148 Muxn ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_out(Muxn_io_out)
  );
  Muxn_148 Muxn_1 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_out(Muxn_1_io_out)
  );
  Muxn_148 Muxn_2 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_in_3(Muxn_2_io_in_3),
    .io_out(Muxn_2_io_out)
  );
  Muxn_148 Muxn_3 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_in_3(Muxn_3_io_in_3),
    .io_out(Muxn_3_io_out)
  );
  Muxn_148 Muxn_4 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_in_3(Muxn_4_io_in_3),
    .io_out(Muxn_4_io_out)
  );
  Muxn_148 Muxn_5 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_in_3(Muxn_5_io_in_3),
    .io_out(Muxn_5_io_out)
  );
  Muxn_148 Muxn_6 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_out(Muxn_6_io_out)
  );
  Muxn_148 Muxn_7 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_out(Muxn_7_io_out)
  );
  Muxn_147 Muxn_8 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_147 Muxn_9 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  Muxn_147 Muxn_10 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_10_io_config),
    .io_in_0(Muxn_10_io_in_0),
    .io_in_1(Muxn_10_io_in_1),
    .io_in_2(Muxn_10_io_in_2),
    .io_in_3(Muxn_10_io_in_3),
    .io_in_4(Muxn_10_io_in_4),
    .io_out(Muxn_10_io_out)
  );
  Muxn_147 Muxn_11 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_11_io_config),
    .io_in_0(Muxn_11_io_in_0),
    .io_in_1(Muxn_11_io_in_1),
    .io_in_2(Muxn_11_io_in_2),
    .io_in_3(Muxn_11_io_in_3),
    .io_in_4(Muxn_11_io_in_4),
    .io_out(Muxn_11_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNE_0 = Muxn_2_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinNE_1 = Muxn_3_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinSE_0 = Muxn_4_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSE_1 = Muxn_5_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSW_0 = Muxn_6_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_ipinSW_1 = Muxn_7_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_otrackW_0 = Muxn_8_io_out; // @[Interconnect.scala 430:21 Interconnect.scala 479:45]
  assign io_otrackN_0 = Muxn_9_io_out; // @[Interconnect.scala 431:21 Interconnect.scala 479:45]
  assign io_otrackE_0 = Muxn_10_io_out; // @[Interconnect.scala 432:21 Interconnect.scala 479:45]
  assign io_otrackS_0 = Muxn_11_io_out; // @[Interconnect.scala 433:21 Interconnect.scala 479:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 464:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 466:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 483:23]
  assign Muxn_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 483:23]
  assign Muxn_1_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 483:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 483:23]
  assign Muxn_3_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 483:23]
  assign Muxn_4_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 483:23]
  assign Muxn_5_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[13:12]; // @[Interconnect.scala 483:23]
  assign Muxn_6_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[15:14]; // @[Interconnect.scala 483:23]
  assign Muxn_7_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[18:16]; // @[Interconnect.scala 483:23]
  assign Muxn_8_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[21:19]; // @[Interconnect.scala 483:23]
  assign Muxn_9_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_config = ConfigMem_io_out_0[24:22]; // @[Interconnect.scala 483:23]
  assign Muxn_10_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_config = ConfigMem_io_out_0[27:25]; // @[Interconnect.scala 483:23]
  assign Muxn_11_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_4 = io_itrackE_0; // @[Interconnect.scala 475:63]
endmodule
module GIB_25(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire  ConfigMem_clock; // @[Interconnect.scala 463:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 463:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 463:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 463:21]
  wire [27:0] ConfigMem_io_out_0; // @[Interconnect.scala 463:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_6_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_7_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_10_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_11_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_out; // @[Interconnect.scala 473:25]
  wire  _T_1 = 10'h3e == io_cfg_addr[11:2]; // @[Interconnect.scala 464:50]
  reg [31:0] _T_12; // @[Interconnect.scala 477:55]
  reg [31:0] _T_14; // @[Interconnect.scala 477:55]
  reg [31:0] _T_16; // @[Interconnect.scala 477:55]
  reg [31:0] _T_18; // @[Interconnect.scala 477:55]
  ConfigMem_90 ConfigMem ( // @[Interconnect.scala 463:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_148 Muxn ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_out(Muxn_io_out)
  );
  Muxn_148 Muxn_1 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_out(Muxn_1_io_out)
  );
  Muxn_148 Muxn_2 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_in_3(Muxn_2_io_in_3),
    .io_out(Muxn_2_io_out)
  );
  Muxn_148 Muxn_3 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_in_3(Muxn_3_io_in_3),
    .io_out(Muxn_3_io_out)
  );
  Muxn_148 Muxn_4 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_in_3(Muxn_4_io_in_3),
    .io_out(Muxn_4_io_out)
  );
  Muxn_148 Muxn_5 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_in_3(Muxn_5_io_in_3),
    .io_out(Muxn_5_io_out)
  );
  Muxn_148 Muxn_6 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_out(Muxn_6_io_out)
  );
  Muxn_148 Muxn_7 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_out(Muxn_7_io_out)
  );
  Muxn_147 Muxn_8 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_147 Muxn_9 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  Muxn_147 Muxn_10 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_10_io_config),
    .io_in_0(Muxn_10_io_in_0),
    .io_in_1(Muxn_10_io_in_1),
    .io_in_2(Muxn_10_io_in_2),
    .io_in_3(Muxn_10_io_in_3),
    .io_in_4(Muxn_10_io_in_4),
    .io_out(Muxn_10_io_out)
  );
  Muxn_147 Muxn_11 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_11_io_config),
    .io_in_0(Muxn_11_io_in_0),
    .io_in_1(Muxn_11_io_in_1),
    .io_in_2(Muxn_11_io_in_2),
    .io_in_3(Muxn_11_io_in_3),
    .io_in_4(Muxn_11_io_in_4),
    .io_out(Muxn_11_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNE_0 = Muxn_2_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinNE_1 = Muxn_3_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinSE_0 = Muxn_4_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSE_1 = Muxn_5_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSW_0 = Muxn_6_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_ipinSW_1 = Muxn_7_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_otrackW_0 = _T_12; // @[Interconnect.scala 430:21 Interconnect.scala 477:45]
  assign io_otrackN_0 = _T_14; // @[Interconnect.scala 431:21 Interconnect.scala 477:45]
  assign io_otrackE_0 = _T_16; // @[Interconnect.scala 432:21 Interconnect.scala 477:45]
  assign io_otrackS_0 = _T_18; // @[Interconnect.scala 433:21 Interconnect.scala 477:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 464:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 466:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 483:23]
  assign Muxn_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 483:23]
  assign Muxn_1_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 483:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 483:23]
  assign Muxn_3_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 483:23]
  assign Muxn_4_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 483:23]
  assign Muxn_5_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[13:12]; // @[Interconnect.scala 483:23]
  assign Muxn_6_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[15:14]; // @[Interconnect.scala 483:23]
  assign Muxn_7_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[18:16]; // @[Interconnect.scala 483:23]
  assign Muxn_8_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[21:19]; // @[Interconnect.scala 483:23]
  assign Muxn_9_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_config = ConfigMem_io_out_0[24:22]; // @[Interconnect.scala 483:23]
  assign Muxn_10_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_config = ConfigMem_io_out_0[27:25]; // @[Interconnect.scala 483:23]
  assign Muxn_11_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_4 = io_itrackE_0; // @[Interconnect.scala 475:63]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_12 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  _T_14 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  _T_16 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  _T_18 = _RAND_3[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_12 <= Muxn_8_io_out;
    _T_14 <= Muxn_9_io_out;
    _T_16 <= Muxn_10_io_out;
    _T_18 <= Muxn_11_io_out;
  end
endmodule
module GIB_26(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
  wire  ConfigMem_clock; // @[Interconnect.scala 463:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 463:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 463:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 463:21]
  wire [14:0] ConfigMem_io_out_0; // @[Interconnect.scala 463:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 473:25]
  wire  Muxn_2_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 473:25]
  wire  Muxn_3_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_6_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_7_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 473:25]
  wire  _T_1 = 10'h3f == io_cfg_addr[11:2]; // @[Interconnect.scala 464:50]
  ConfigMem_89 ConfigMem ( // @[Interconnect.scala 463:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_145 Muxn ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_out(Muxn_io_out)
  );
  Muxn_145 Muxn_1 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_out(Muxn_1_io_out)
  );
  Muxn Muxn_2 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_out(Muxn_2_io_out)
  );
  Muxn Muxn_3 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_out(Muxn_3_io_out)
  );
  Muxn_145 Muxn_4 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_out(Muxn_4_io_out)
  );
  Muxn_148 Muxn_5 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_in_3(Muxn_5_io_in_3),
    .io_out(Muxn_5_io_out)
  );
  Muxn_147 Muxn_6 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_in_4(Muxn_6_io_in_4),
    .io_out(Muxn_6_io_out)
  );
  Muxn_148 Muxn_7 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_out(Muxn_7_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinSW_0 = Muxn_2_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_ipinSW_1 = Muxn_3_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_otrackW_0 = Muxn_4_io_out; // @[Interconnect.scala 430:21 Interconnect.scala 479:45]
  assign io_otrackN_0 = Muxn_5_io_out; // @[Interconnect.scala 431:21 Interconnect.scala 479:45]
  assign io_otrackS_0 = Muxn_7_io_out; // @[Interconnect.scala 433:21 Interconnect.scala 479:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 464:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 466:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 483:23]
  assign Muxn_io_in_0 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_1 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_2 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 483:23]
  assign Muxn_1_io_in_0 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_1 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_2 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[4]; // @[Interconnect.scala 483:23]
  assign Muxn_2_io_in_0 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_1 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[5]; // @[Interconnect.scala 483:23]
  assign Muxn_3_io_in_0 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_1 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 483:23]
  assign Muxn_4_io_in_0 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_1 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_2 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 483:23]
  assign Muxn_5_io_in_0 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_1 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_2 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[12:10]; // @[Interconnect.scala 483:23]
  assign Muxn_6_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[14:13]; // @[Interconnect.scala 483:23]
  assign Muxn_7_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_1 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_3 = 32'h0; // @[Interconnect.scala 475:63]
endmodule
module GIB_27(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire  ConfigMem_clock; // @[Interconnect.scala 463:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 463:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 463:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 463:21]
  wire [14:0] ConfigMem_io_out_0; // @[Interconnect.scala 463:21]
  wire  Muxn_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 473:25]
  wire  Muxn_1_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_4_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_6_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_7_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 473:25]
  wire  _T_1 = 10'h49 == io_cfg_addr[11:2]; // @[Interconnect.scala 464:50]
  reg [31:0] _T_10; // @[Interconnect.scala 477:55]
  reg [31:0] _T_12; // @[Interconnect.scala 477:55]
  reg [31:0] _T_14; // @[Interconnect.scala 477:55]
  ConfigMem_89 ConfigMem ( // @[Interconnect.scala 463:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn Muxn ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_out(Muxn_io_out)
  );
  Muxn Muxn_1 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_out(Muxn_1_io_out)
  );
  Muxn_145 Muxn_2 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_out(Muxn_2_io_out)
  );
  Muxn_145 Muxn_3 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_out(Muxn_3_io_out)
  );
  Muxn_147 Muxn_4 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_in_3(Muxn_4_io_in_3),
    .io_in_4(Muxn_4_io_in_4),
    .io_out(Muxn_4_io_out)
  );
  Muxn_148 Muxn_5 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_in_3(Muxn_5_io_in_3),
    .io_out(Muxn_5_io_out)
  );
  Muxn_145 Muxn_6 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_out(Muxn_6_io_out)
  );
  Muxn_148 Muxn_7 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_out(Muxn_7_io_out)
  );
  assign io_ipinNE_0 = Muxn_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinNE_1 = Muxn_1_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinSE_0 = Muxn_2_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSE_1 = Muxn_3_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_otrackN_0 = _T_10; // @[Interconnect.scala 431:21 Interconnect.scala 477:45]
  assign io_otrackE_0 = _T_12; // @[Interconnect.scala 432:21 Interconnect.scala 477:45]
  assign io_otrackS_0 = _T_14; // @[Interconnect.scala 433:21 Interconnect.scala 477:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 464:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 466:21]
  assign Muxn_io_config = ConfigMem_io_out_0[0]; // @[Interconnect.scala 483:23]
  assign Muxn_io_in_0 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_1 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[1]; // @[Interconnect.scala 483:23]
  assign Muxn_1_io_in_0 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_1 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 483:23]
  assign Muxn_2_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_1 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 483:23]
  assign Muxn_3_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_1 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[8:6]; // @[Interconnect.scala 483:23]
  assign Muxn_4_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[10:9]; // @[Interconnect.scala 483:23]
  assign Muxn_5_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_1 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[12:11]; // @[Interconnect.scala 483:23]
  assign Muxn_6_io_in_0 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_1 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_2 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[14:13]; // @[Interconnect.scala 483:23]
  assign Muxn_7_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_1 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_10 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  _T_12 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  _T_14 = _RAND_2[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_10 <= Muxn_5_io_out;
    _T_12 <= Muxn_6_io_out;
    _T_14 <= Muxn_7_io_out;
  end
endmodule
module GIB_28(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
  wire  ConfigMem_clock; // @[Interconnect.scala 463:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 463:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 463:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 463:21]
  wire [27:0] ConfigMem_io_out_0; // @[Interconnect.scala 463:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_6_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_7_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_10_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_11_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_out; // @[Interconnect.scala 473:25]
  wire  _T_1 = 10'h4a == io_cfg_addr[11:2]; // @[Interconnect.scala 464:50]
  ConfigMem_90 ConfigMem ( // @[Interconnect.scala 463:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_148 Muxn ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_out(Muxn_io_out)
  );
  Muxn_148 Muxn_1 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_out(Muxn_1_io_out)
  );
  Muxn_148 Muxn_2 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_in_3(Muxn_2_io_in_3),
    .io_out(Muxn_2_io_out)
  );
  Muxn_148 Muxn_3 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_in_3(Muxn_3_io_in_3),
    .io_out(Muxn_3_io_out)
  );
  Muxn_148 Muxn_4 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_in_3(Muxn_4_io_in_3),
    .io_out(Muxn_4_io_out)
  );
  Muxn_148 Muxn_5 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_in_3(Muxn_5_io_in_3),
    .io_out(Muxn_5_io_out)
  );
  Muxn_148 Muxn_6 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_out(Muxn_6_io_out)
  );
  Muxn_148 Muxn_7 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_out(Muxn_7_io_out)
  );
  Muxn_147 Muxn_8 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_147 Muxn_9 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  Muxn_147 Muxn_10 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_10_io_config),
    .io_in_0(Muxn_10_io_in_0),
    .io_in_1(Muxn_10_io_in_1),
    .io_in_2(Muxn_10_io_in_2),
    .io_in_3(Muxn_10_io_in_3),
    .io_in_4(Muxn_10_io_in_4),
    .io_out(Muxn_10_io_out)
  );
  Muxn_147 Muxn_11 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_11_io_config),
    .io_in_0(Muxn_11_io_in_0),
    .io_in_1(Muxn_11_io_in_1),
    .io_in_2(Muxn_11_io_in_2),
    .io_in_3(Muxn_11_io_in_3),
    .io_in_4(Muxn_11_io_in_4),
    .io_out(Muxn_11_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNE_0 = Muxn_2_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinNE_1 = Muxn_3_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinSE_0 = Muxn_4_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSE_1 = Muxn_5_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSW_0 = Muxn_6_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_ipinSW_1 = Muxn_7_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_otrackW_0 = Muxn_8_io_out; // @[Interconnect.scala 430:21 Interconnect.scala 479:45]
  assign io_otrackN_0 = Muxn_9_io_out; // @[Interconnect.scala 431:21 Interconnect.scala 479:45]
  assign io_otrackE_0 = Muxn_10_io_out; // @[Interconnect.scala 432:21 Interconnect.scala 479:45]
  assign io_otrackS_0 = Muxn_11_io_out; // @[Interconnect.scala 433:21 Interconnect.scala 479:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 464:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 466:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 483:23]
  assign Muxn_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 483:23]
  assign Muxn_1_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 483:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 483:23]
  assign Muxn_3_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 483:23]
  assign Muxn_4_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 483:23]
  assign Muxn_5_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[13:12]; // @[Interconnect.scala 483:23]
  assign Muxn_6_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[15:14]; // @[Interconnect.scala 483:23]
  assign Muxn_7_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[18:16]; // @[Interconnect.scala 483:23]
  assign Muxn_8_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[21:19]; // @[Interconnect.scala 483:23]
  assign Muxn_9_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_config = ConfigMem_io_out_0[24:22]; // @[Interconnect.scala 483:23]
  assign Muxn_10_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_config = ConfigMem_io_out_0[27:25]; // @[Interconnect.scala 483:23]
  assign Muxn_11_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_4 = io_itrackE_0; // @[Interconnect.scala 475:63]
endmodule
module GIB_29(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire  ConfigMem_clock; // @[Interconnect.scala 463:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 463:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 463:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 463:21]
  wire [27:0] ConfigMem_io_out_0; // @[Interconnect.scala 463:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_6_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_7_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_10_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_11_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_out; // @[Interconnect.scala 473:25]
  wire  _T_1 = 10'h4b == io_cfg_addr[11:2]; // @[Interconnect.scala 464:50]
  reg [31:0] _T_12; // @[Interconnect.scala 477:55]
  reg [31:0] _T_14; // @[Interconnect.scala 477:55]
  reg [31:0] _T_16; // @[Interconnect.scala 477:55]
  reg [31:0] _T_18; // @[Interconnect.scala 477:55]
  ConfigMem_90 ConfigMem ( // @[Interconnect.scala 463:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_148 Muxn ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_out(Muxn_io_out)
  );
  Muxn_148 Muxn_1 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_out(Muxn_1_io_out)
  );
  Muxn_148 Muxn_2 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_in_3(Muxn_2_io_in_3),
    .io_out(Muxn_2_io_out)
  );
  Muxn_148 Muxn_3 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_in_3(Muxn_3_io_in_3),
    .io_out(Muxn_3_io_out)
  );
  Muxn_148 Muxn_4 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_in_3(Muxn_4_io_in_3),
    .io_out(Muxn_4_io_out)
  );
  Muxn_148 Muxn_5 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_in_3(Muxn_5_io_in_3),
    .io_out(Muxn_5_io_out)
  );
  Muxn_148 Muxn_6 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_out(Muxn_6_io_out)
  );
  Muxn_148 Muxn_7 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_out(Muxn_7_io_out)
  );
  Muxn_147 Muxn_8 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_147 Muxn_9 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  Muxn_147 Muxn_10 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_10_io_config),
    .io_in_0(Muxn_10_io_in_0),
    .io_in_1(Muxn_10_io_in_1),
    .io_in_2(Muxn_10_io_in_2),
    .io_in_3(Muxn_10_io_in_3),
    .io_in_4(Muxn_10_io_in_4),
    .io_out(Muxn_10_io_out)
  );
  Muxn_147 Muxn_11 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_11_io_config),
    .io_in_0(Muxn_11_io_in_0),
    .io_in_1(Muxn_11_io_in_1),
    .io_in_2(Muxn_11_io_in_2),
    .io_in_3(Muxn_11_io_in_3),
    .io_in_4(Muxn_11_io_in_4),
    .io_out(Muxn_11_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNE_0 = Muxn_2_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinNE_1 = Muxn_3_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinSE_0 = Muxn_4_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSE_1 = Muxn_5_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSW_0 = Muxn_6_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_ipinSW_1 = Muxn_7_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_otrackW_0 = _T_12; // @[Interconnect.scala 430:21 Interconnect.scala 477:45]
  assign io_otrackN_0 = _T_14; // @[Interconnect.scala 431:21 Interconnect.scala 477:45]
  assign io_otrackE_0 = _T_16; // @[Interconnect.scala 432:21 Interconnect.scala 477:45]
  assign io_otrackS_0 = _T_18; // @[Interconnect.scala 433:21 Interconnect.scala 477:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 464:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 466:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 483:23]
  assign Muxn_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 483:23]
  assign Muxn_1_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 483:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 483:23]
  assign Muxn_3_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 483:23]
  assign Muxn_4_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 483:23]
  assign Muxn_5_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[13:12]; // @[Interconnect.scala 483:23]
  assign Muxn_6_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[15:14]; // @[Interconnect.scala 483:23]
  assign Muxn_7_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[18:16]; // @[Interconnect.scala 483:23]
  assign Muxn_8_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[21:19]; // @[Interconnect.scala 483:23]
  assign Muxn_9_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_config = ConfigMem_io_out_0[24:22]; // @[Interconnect.scala 483:23]
  assign Muxn_10_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_config = ConfigMem_io_out_0[27:25]; // @[Interconnect.scala 483:23]
  assign Muxn_11_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_4 = io_itrackE_0; // @[Interconnect.scala 475:63]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_12 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  _T_14 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  _T_16 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  _T_18 = _RAND_3[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_12 <= Muxn_8_io_out;
    _T_14 <= Muxn_9_io_out;
    _T_16 <= Muxn_10_io_out;
    _T_18 <= Muxn_11_io_out;
  end
endmodule
module GIB_30(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
  wire  ConfigMem_clock; // @[Interconnect.scala 463:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 463:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 463:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 463:21]
  wire [27:0] ConfigMem_io_out_0; // @[Interconnect.scala 463:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_6_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_7_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_10_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_11_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_out; // @[Interconnect.scala 473:25]
  wire  _T_1 = 10'h4c == io_cfg_addr[11:2]; // @[Interconnect.scala 464:50]
  ConfigMem_90 ConfigMem ( // @[Interconnect.scala 463:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_148 Muxn ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_out(Muxn_io_out)
  );
  Muxn_148 Muxn_1 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_out(Muxn_1_io_out)
  );
  Muxn_148 Muxn_2 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_in_3(Muxn_2_io_in_3),
    .io_out(Muxn_2_io_out)
  );
  Muxn_148 Muxn_3 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_in_3(Muxn_3_io_in_3),
    .io_out(Muxn_3_io_out)
  );
  Muxn_148 Muxn_4 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_in_3(Muxn_4_io_in_3),
    .io_out(Muxn_4_io_out)
  );
  Muxn_148 Muxn_5 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_in_3(Muxn_5_io_in_3),
    .io_out(Muxn_5_io_out)
  );
  Muxn_148 Muxn_6 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_out(Muxn_6_io_out)
  );
  Muxn_148 Muxn_7 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_out(Muxn_7_io_out)
  );
  Muxn_147 Muxn_8 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_147 Muxn_9 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  Muxn_147 Muxn_10 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_10_io_config),
    .io_in_0(Muxn_10_io_in_0),
    .io_in_1(Muxn_10_io_in_1),
    .io_in_2(Muxn_10_io_in_2),
    .io_in_3(Muxn_10_io_in_3),
    .io_in_4(Muxn_10_io_in_4),
    .io_out(Muxn_10_io_out)
  );
  Muxn_147 Muxn_11 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_11_io_config),
    .io_in_0(Muxn_11_io_in_0),
    .io_in_1(Muxn_11_io_in_1),
    .io_in_2(Muxn_11_io_in_2),
    .io_in_3(Muxn_11_io_in_3),
    .io_in_4(Muxn_11_io_in_4),
    .io_out(Muxn_11_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNE_0 = Muxn_2_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinNE_1 = Muxn_3_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinSE_0 = Muxn_4_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSE_1 = Muxn_5_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSW_0 = Muxn_6_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_ipinSW_1 = Muxn_7_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_otrackW_0 = Muxn_8_io_out; // @[Interconnect.scala 430:21 Interconnect.scala 479:45]
  assign io_otrackN_0 = Muxn_9_io_out; // @[Interconnect.scala 431:21 Interconnect.scala 479:45]
  assign io_otrackE_0 = Muxn_10_io_out; // @[Interconnect.scala 432:21 Interconnect.scala 479:45]
  assign io_otrackS_0 = Muxn_11_io_out; // @[Interconnect.scala 433:21 Interconnect.scala 479:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 464:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 466:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 483:23]
  assign Muxn_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 483:23]
  assign Muxn_1_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 483:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 483:23]
  assign Muxn_3_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 483:23]
  assign Muxn_4_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 483:23]
  assign Muxn_5_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[13:12]; // @[Interconnect.scala 483:23]
  assign Muxn_6_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[15:14]; // @[Interconnect.scala 483:23]
  assign Muxn_7_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[18:16]; // @[Interconnect.scala 483:23]
  assign Muxn_8_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[21:19]; // @[Interconnect.scala 483:23]
  assign Muxn_9_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_config = ConfigMem_io_out_0[24:22]; // @[Interconnect.scala 483:23]
  assign Muxn_10_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_config = ConfigMem_io_out_0[27:25]; // @[Interconnect.scala 483:23]
  assign Muxn_11_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_4 = io_itrackE_0; // @[Interconnect.scala 475:63]
endmodule
module GIB_31(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire  ConfigMem_clock; // @[Interconnect.scala 463:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 463:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 463:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 463:21]
  wire [27:0] ConfigMem_io_out_0; // @[Interconnect.scala 463:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_6_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_7_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_10_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_11_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_out; // @[Interconnect.scala 473:25]
  wire  _T_1 = 10'h4d == io_cfg_addr[11:2]; // @[Interconnect.scala 464:50]
  reg [31:0] _T_12; // @[Interconnect.scala 477:55]
  reg [31:0] _T_14; // @[Interconnect.scala 477:55]
  reg [31:0] _T_16; // @[Interconnect.scala 477:55]
  reg [31:0] _T_18; // @[Interconnect.scala 477:55]
  ConfigMem_90 ConfigMem ( // @[Interconnect.scala 463:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_148 Muxn ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_out(Muxn_io_out)
  );
  Muxn_148 Muxn_1 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_out(Muxn_1_io_out)
  );
  Muxn_148 Muxn_2 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_in_3(Muxn_2_io_in_3),
    .io_out(Muxn_2_io_out)
  );
  Muxn_148 Muxn_3 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_in_3(Muxn_3_io_in_3),
    .io_out(Muxn_3_io_out)
  );
  Muxn_148 Muxn_4 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_in_3(Muxn_4_io_in_3),
    .io_out(Muxn_4_io_out)
  );
  Muxn_148 Muxn_5 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_in_3(Muxn_5_io_in_3),
    .io_out(Muxn_5_io_out)
  );
  Muxn_148 Muxn_6 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_out(Muxn_6_io_out)
  );
  Muxn_148 Muxn_7 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_out(Muxn_7_io_out)
  );
  Muxn_147 Muxn_8 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_147 Muxn_9 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  Muxn_147 Muxn_10 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_10_io_config),
    .io_in_0(Muxn_10_io_in_0),
    .io_in_1(Muxn_10_io_in_1),
    .io_in_2(Muxn_10_io_in_2),
    .io_in_3(Muxn_10_io_in_3),
    .io_in_4(Muxn_10_io_in_4),
    .io_out(Muxn_10_io_out)
  );
  Muxn_147 Muxn_11 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_11_io_config),
    .io_in_0(Muxn_11_io_in_0),
    .io_in_1(Muxn_11_io_in_1),
    .io_in_2(Muxn_11_io_in_2),
    .io_in_3(Muxn_11_io_in_3),
    .io_in_4(Muxn_11_io_in_4),
    .io_out(Muxn_11_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNE_0 = Muxn_2_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinNE_1 = Muxn_3_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinSE_0 = Muxn_4_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSE_1 = Muxn_5_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSW_0 = Muxn_6_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_ipinSW_1 = Muxn_7_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_otrackW_0 = _T_12; // @[Interconnect.scala 430:21 Interconnect.scala 477:45]
  assign io_otrackN_0 = _T_14; // @[Interconnect.scala 431:21 Interconnect.scala 477:45]
  assign io_otrackE_0 = _T_16; // @[Interconnect.scala 432:21 Interconnect.scala 477:45]
  assign io_otrackS_0 = _T_18; // @[Interconnect.scala 433:21 Interconnect.scala 477:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 464:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 466:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 483:23]
  assign Muxn_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 483:23]
  assign Muxn_1_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 483:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 483:23]
  assign Muxn_3_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 483:23]
  assign Muxn_4_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 483:23]
  assign Muxn_5_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[13:12]; // @[Interconnect.scala 483:23]
  assign Muxn_6_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[15:14]; // @[Interconnect.scala 483:23]
  assign Muxn_7_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[18:16]; // @[Interconnect.scala 483:23]
  assign Muxn_8_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[21:19]; // @[Interconnect.scala 483:23]
  assign Muxn_9_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_config = ConfigMem_io_out_0[24:22]; // @[Interconnect.scala 483:23]
  assign Muxn_10_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_config = ConfigMem_io_out_0[27:25]; // @[Interconnect.scala 483:23]
  assign Muxn_11_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_4 = io_itrackE_0; // @[Interconnect.scala 475:63]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_12 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  _T_14 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  _T_16 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  _T_18 = _RAND_3[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_12 <= Muxn_8_io_out;
    _T_14 <= Muxn_9_io_out;
    _T_16 <= Muxn_10_io_out;
    _T_18 <= Muxn_11_io_out;
  end
endmodule
module GIB_32(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
  wire  ConfigMem_clock; // @[Interconnect.scala 463:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 463:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 463:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 463:21]
  wire [27:0] ConfigMem_io_out_0; // @[Interconnect.scala 463:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_6_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_7_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_10_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_11_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_out; // @[Interconnect.scala 473:25]
  wire  _T_1 = 10'h4e == io_cfg_addr[11:2]; // @[Interconnect.scala 464:50]
  ConfigMem_90 ConfigMem ( // @[Interconnect.scala 463:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_148 Muxn ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_out(Muxn_io_out)
  );
  Muxn_148 Muxn_1 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_out(Muxn_1_io_out)
  );
  Muxn_148 Muxn_2 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_in_3(Muxn_2_io_in_3),
    .io_out(Muxn_2_io_out)
  );
  Muxn_148 Muxn_3 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_in_3(Muxn_3_io_in_3),
    .io_out(Muxn_3_io_out)
  );
  Muxn_148 Muxn_4 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_in_3(Muxn_4_io_in_3),
    .io_out(Muxn_4_io_out)
  );
  Muxn_148 Muxn_5 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_in_3(Muxn_5_io_in_3),
    .io_out(Muxn_5_io_out)
  );
  Muxn_148 Muxn_6 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_out(Muxn_6_io_out)
  );
  Muxn_148 Muxn_7 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_out(Muxn_7_io_out)
  );
  Muxn_147 Muxn_8 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_147 Muxn_9 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  Muxn_147 Muxn_10 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_10_io_config),
    .io_in_0(Muxn_10_io_in_0),
    .io_in_1(Muxn_10_io_in_1),
    .io_in_2(Muxn_10_io_in_2),
    .io_in_3(Muxn_10_io_in_3),
    .io_in_4(Muxn_10_io_in_4),
    .io_out(Muxn_10_io_out)
  );
  Muxn_147 Muxn_11 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_11_io_config),
    .io_in_0(Muxn_11_io_in_0),
    .io_in_1(Muxn_11_io_in_1),
    .io_in_2(Muxn_11_io_in_2),
    .io_in_3(Muxn_11_io_in_3),
    .io_in_4(Muxn_11_io_in_4),
    .io_out(Muxn_11_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNE_0 = Muxn_2_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinNE_1 = Muxn_3_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinSE_0 = Muxn_4_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSE_1 = Muxn_5_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSW_0 = Muxn_6_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_ipinSW_1 = Muxn_7_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_otrackW_0 = Muxn_8_io_out; // @[Interconnect.scala 430:21 Interconnect.scala 479:45]
  assign io_otrackN_0 = Muxn_9_io_out; // @[Interconnect.scala 431:21 Interconnect.scala 479:45]
  assign io_otrackE_0 = Muxn_10_io_out; // @[Interconnect.scala 432:21 Interconnect.scala 479:45]
  assign io_otrackS_0 = Muxn_11_io_out; // @[Interconnect.scala 433:21 Interconnect.scala 479:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 464:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 466:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 483:23]
  assign Muxn_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 483:23]
  assign Muxn_1_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 483:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 483:23]
  assign Muxn_3_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 483:23]
  assign Muxn_4_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 483:23]
  assign Muxn_5_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[13:12]; // @[Interconnect.scala 483:23]
  assign Muxn_6_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[15:14]; // @[Interconnect.scala 483:23]
  assign Muxn_7_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[18:16]; // @[Interconnect.scala 483:23]
  assign Muxn_8_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[21:19]; // @[Interconnect.scala 483:23]
  assign Muxn_9_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_config = ConfigMem_io_out_0[24:22]; // @[Interconnect.scala 483:23]
  assign Muxn_10_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_config = ConfigMem_io_out_0[27:25]; // @[Interconnect.scala 483:23]
  assign Muxn_11_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_4 = io_itrackE_0; // @[Interconnect.scala 475:63]
endmodule
module GIB_33(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire  ConfigMem_clock; // @[Interconnect.scala 463:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 463:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 463:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 463:21]
  wire [27:0] ConfigMem_io_out_0; // @[Interconnect.scala 463:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_6_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_7_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_10_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_11_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_out; // @[Interconnect.scala 473:25]
  wire  _T_1 = 10'h4f == io_cfg_addr[11:2]; // @[Interconnect.scala 464:50]
  reg [31:0] _T_12; // @[Interconnect.scala 477:55]
  reg [31:0] _T_14; // @[Interconnect.scala 477:55]
  reg [31:0] _T_16; // @[Interconnect.scala 477:55]
  reg [31:0] _T_18; // @[Interconnect.scala 477:55]
  ConfigMem_90 ConfigMem ( // @[Interconnect.scala 463:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_148 Muxn ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_out(Muxn_io_out)
  );
  Muxn_148 Muxn_1 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_out(Muxn_1_io_out)
  );
  Muxn_148 Muxn_2 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_in_3(Muxn_2_io_in_3),
    .io_out(Muxn_2_io_out)
  );
  Muxn_148 Muxn_3 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_in_3(Muxn_3_io_in_3),
    .io_out(Muxn_3_io_out)
  );
  Muxn_148 Muxn_4 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_in_3(Muxn_4_io_in_3),
    .io_out(Muxn_4_io_out)
  );
  Muxn_148 Muxn_5 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_in_3(Muxn_5_io_in_3),
    .io_out(Muxn_5_io_out)
  );
  Muxn_148 Muxn_6 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_out(Muxn_6_io_out)
  );
  Muxn_148 Muxn_7 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_out(Muxn_7_io_out)
  );
  Muxn_147 Muxn_8 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_147 Muxn_9 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  Muxn_147 Muxn_10 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_10_io_config),
    .io_in_0(Muxn_10_io_in_0),
    .io_in_1(Muxn_10_io_in_1),
    .io_in_2(Muxn_10_io_in_2),
    .io_in_3(Muxn_10_io_in_3),
    .io_in_4(Muxn_10_io_in_4),
    .io_out(Muxn_10_io_out)
  );
  Muxn_147 Muxn_11 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_11_io_config),
    .io_in_0(Muxn_11_io_in_0),
    .io_in_1(Muxn_11_io_in_1),
    .io_in_2(Muxn_11_io_in_2),
    .io_in_3(Muxn_11_io_in_3),
    .io_in_4(Muxn_11_io_in_4),
    .io_out(Muxn_11_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNE_0 = Muxn_2_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinNE_1 = Muxn_3_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinSE_0 = Muxn_4_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSE_1 = Muxn_5_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSW_0 = Muxn_6_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_ipinSW_1 = Muxn_7_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_otrackW_0 = _T_12; // @[Interconnect.scala 430:21 Interconnect.scala 477:45]
  assign io_otrackN_0 = _T_14; // @[Interconnect.scala 431:21 Interconnect.scala 477:45]
  assign io_otrackE_0 = _T_16; // @[Interconnect.scala 432:21 Interconnect.scala 477:45]
  assign io_otrackS_0 = _T_18; // @[Interconnect.scala 433:21 Interconnect.scala 477:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 464:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 466:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 483:23]
  assign Muxn_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 483:23]
  assign Muxn_1_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 483:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 483:23]
  assign Muxn_3_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 483:23]
  assign Muxn_4_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 483:23]
  assign Muxn_5_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[13:12]; // @[Interconnect.scala 483:23]
  assign Muxn_6_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[15:14]; // @[Interconnect.scala 483:23]
  assign Muxn_7_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[18:16]; // @[Interconnect.scala 483:23]
  assign Muxn_8_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[21:19]; // @[Interconnect.scala 483:23]
  assign Muxn_9_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_config = ConfigMem_io_out_0[24:22]; // @[Interconnect.scala 483:23]
  assign Muxn_10_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_config = ConfigMem_io_out_0[27:25]; // @[Interconnect.scala 483:23]
  assign Muxn_11_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_4 = io_itrackE_0; // @[Interconnect.scala 475:63]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_12 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  _T_14 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  _T_16 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  _T_18 = _RAND_3[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_12 <= Muxn_8_io_out;
    _T_14 <= Muxn_9_io_out;
    _T_16 <= Muxn_10_io_out;
    _T_18 <= Muxn_11_io_out;
  end
endmodule
module GIB_34(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
  wire  ConfigMem_clock; // @[Interconnect.scala 463:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 463:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 463:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 463:21]
  wire [27:0] ConfigMem_io_out_0; // @[Interconnect.scala 463:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_6_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_7_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_10_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_11_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_out; // @[Interconnect.scala 473:25]
  wire  _T_1 = 10'h50 == io_cfg_addr[11:2]; // @[Interconnect.scala 464:50]
  ConfigMem_90 ConfigMem ( // @[Interconnect.scala 463:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_148 Muxn ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_out(Muxn_io_out)
  );
  Muxn_148 Muxn_1 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_out(Muxn_1_io_out)
  );
  Muxn_148 Muxn_2 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_in_3(Muxn_2_io_in_3),
    .io_out(Muxn_2_io_out)
  );
  Muxn_148 Muxn_3 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_in_3(Muxn_3_io_in_3),
    .io_out(Muxn_3_io_out)
  );
  Muxn_148 Muxn_4 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_in_3(Muxn_4_io_in_3),
    .io_out(Muxn_4_io_out)
  );
  Muxn_148 Muxn_5 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_in_3(Muxn_5_io_in_3),
    .io_out(Muxn_5_io_out)
  );
  Muxn_148 Muxn_6 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_out(Muxn_6_io_out)
  );
  Muxn_148 Muxn_7 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_out(Muxn_7_io_out)
  );
  Muxn_147 Muxn_8 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_147 Muxn_9 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  Muxn_147 Muxn_10 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_10_io_config),
    .io_in_0(Muxn_10_io_in_0),
    .io_in_1(Muxn_10_io_in_1),
    .io_in_2(Muxn_10_io_in_2),
    .io_in_3(Muxn_10_io_in_3),
    .io_in_4(Muxn_10_io_in_4),
    .io_out(Muxn_10_io_out)
  );
  Muxn_147 Muxn_11 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_11_io_config),
    .io_in_0(Muxn_11_io_in_0),
    .io_in_1(Muxn_11_io_in_1),
    .io_in_2(Muxn_11_io_in_2),
    .io_in_3(Muxn_11_io_in_3),
    .io_in_4(Muxn_11_io_in_4),
    .io_out(Muxn_11_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNE_0 = Muxn_2_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinNE_1 = Muxn_3_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinSE_0 = Muxn_4_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSE_1 = Muxn_5_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSW_0 = Muxn_6_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_ipinSW_1 = Muxn_7_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_otrackW_0 = Muxn_8_io_out; // @[Interconnect.scala 430:21 Interconnect.scala 479:45]
  assign io_otrackN_0 = Muxn_9_io_out; // @[Interconnect.scala 431:21 Interconnect.scala 479:45]
  assign io_otrackE_0 = Muxn_10_io_out; // @[Interconnect.scala 432:21 Interconnect.scala 479:45]
  assign io_otrackS_0 = Muxn_11_io_out; // @[Interconnect.scala 433:21 Interconnect.scala 479:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 464:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 466:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 483:23]
  assign Muxn_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 483:23]
  assign Muxn_1_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 483:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 483:23]
  assign Muxn_3_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 483:23]
  assign Muxn_4_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 483:23]
  assign Muxn_5_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[13:12]; // @[Interconnect.scala 483:23]
  assign Muxn_6_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[15:14]; // @[Interconnect.scala 483:23]
  assign Muxn_7_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[18:16]; // @[Interconnect.scala 483:23]
  assign Muxn_8_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[21:19]; // @[Interconnect.scala 483:23]
  assign Muxn_9_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_config = ConfigMem_io_out_0[24:22]; // @[Interconnect.scala 483:23]
  assign Muxn_10_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_config = ConfigMem_io_out_0[27:25]; // @[Interconnect.scala 483:23]
  assign Muxn_11_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_4 = io_itrackE_0; // @[Interconnect.scala 475:63]
endmodule
module GIB_35(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire  ConfigMem_clock; // @[Interconnect.scala 463:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 463:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 463:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 463:21]
  wire [14:0] ConfigMem_io_out_0; // @[Interconnect.scala 463:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 473:25]
  wire  Muxn_2_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 473:25]
  wire  Muxn_3_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_6_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_7_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 473:25]
  wire  _T_1 = 10'h51 == io_cfg_addr[11:2]; // @[Interconnect.scala 464:50]
  reg [31:0] _T_8; // @[Interconnect.scala 477:55]
  reg [31:0] _T_10; // @[Interconnect.scala 477:55]
  reg [31:0] _T_14; // @[Interconnect.scala 477:55]
  ConfigMem_89 ConfigMem ( // @[Interconnect.scala 463:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_145 Muxn ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_out(Muxn_io_out)
  );
  Muxn_145 Muxn_1 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_out(Muxn_1_io_out)
  );
  Muxn Muxn_2 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_out(Muxn_2_io_out)
  );
  Muxn Muxn_3 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_out(Muxn_3_io_out)
  );
  Muxn_145 Muxn_4 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_out(Muxn_4_io_out)
  );
  Muxn_148 Muxn_5 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_in_3(Muxn_5_io_in_3),
    .io_out(Muxn_5_io_out)
  );
  Muxn_147 Muxn_6 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_in_4(Muxn_6_io_in_4),
    .io_out(Muxn_6_io_out)
  );
  Muxn_148 Muxn_7 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_out(Muxn_7_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinSW_0 = Muxn_2_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_ipinSW_1 = Muxn_3_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_otrackW_0 = _T_8; // @[Interconnect.scala 430:21 Interconnect.scala 477:45]
  assign io_otrackN_0 = _T_10; // @[Interconnect.scala 431:21 Interconnect.scala 477:45]
  assign io_otrackS_0 = _T_14; // @[Interconnect.scala 433:21 Interconnect.scala 477:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 464:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 466:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 483:23]
  assign Muxn_io_in_0 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_1 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_2 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 483:23]
  assign Muxn_1_io_in_0 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_1 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_2 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[4]; // @[Interconnect.scala 483:23]
  assign Muxn_2_io_in_0 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_1 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[5]; // @[Interconnect.scala 483:23]
  assign Muxn_3_io_in_0 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_1 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 483:23]
  assign Muxn_4_io_in_0 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_1 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_2 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 483:23]
  assign Muxn_5_io_in_0 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_1 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_2 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[12:10]; // @[Interconnect.scala 483:23]
  assign Muxn_6_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[14:13]; // @[Interconnect.scala 483:23]
  assign Muxn_7_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_1 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_3 = 32'h0; // @[Interconnect.scala 475:63]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_8 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  _T_10 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  _T_14 = _RAND_2[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_8 <= Muxn_4_io_out;
    _T_10 <= Muxn_5_io_out;
    _T_14 <= Muxn_7_io_out;
  end
endmodule
module GIB_36(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
  wire  ConfigMem_clock; // @[Interconnect.scala 463:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 463:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 463:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 463:21]
  wire [14:0] ConfigMem_io_out_0; // @[Interconnect.scala 463:21]
  wire  Muxn_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 473:25]
  wire  Muxn_1_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_4_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_6_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_7_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 473:25]
  wire  _T_1 = 10'h5b == io_cfg_addr[11:2]; // @[Interconnect.scala 464:50]
  ConfigMem_89 ConfigMem ( // @[Interconnect.scala 463:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn Muxn ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_out(Muxn_io_out)
  );
  Muxn Muxn_1 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_out(Muxn_1_io_out)
  );
  Muxn_145 Muxn_2 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_out(Muxn_2_io_out)
  );
  Muxn_145 Muxn_3 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_out(Muxn_3_io_out)
  );
  Muxn_147 Muxn_4 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_in_3(Muxn_4_io_in_3),
    .io_in_4(Muxn_4_io_in_4),
    .io_out(Muxn_4_io_out)
  );
  Muxn_148 Muxn_5 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_in_3(Muxn_5_io_in_3),
    .io_out(Muxn_5_io_out)
  );
  Muxn_145 Muxn_6 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_out(Muxn_6_io_out)
  );
  Muxn_148 Muxn_7 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_out(Muxn_7_io_out)
  );
  assign io_ipinNE_0 = Muxn_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinNE_1 = Muxn_1_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinSE_0 = Muxn_2_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSE_1 = Muxn_3_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_otrackN_0 = Muxn_5_io_out; // @[Interconnect.scala 431:21 Interconnect.scala 479:45]
  assign io_otrackE_0 = Muxn_6_io_out; // @[Interconnect.scala 432:21 Interconnect.scala 479:45]
  assign io_otrackS_0 = Muxn_7_io_out; // @[Interconnect.scala 433:21 Interconnect.scala 479:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 464:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 466:21]
  assign Muxn_io_config = ConfigMem_io_out_0[0]; // @[Interconnect.scala 483:23]
  assign Muxn_io_in_0 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_1 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[1]; // @[Interconnect.scala 483:23]
  assign Muxn_1_io_in_0 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_1 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 483:23]
  assign Muxn_2_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_1 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 483:23]
  assign Muxn_3_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_1 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[8:6]; // @[Interconnect.scala 483:23]
  assign Muxn_4_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[10:9]; // @[Interconnect.scala 483:23]
  assign Muxn_5_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_1 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[12:11]; // @[Interconnect.scala 483:23]
  assign Muxn_6_io_in_0 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_1 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_2 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[14:13]; // @[Interconnect.scala 483:23]
  assign Muxn_7_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_1 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
endmodule
module GIB_37(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire  ConfigMem_clock; // @[Interconnect.scala 463:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 463:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 463:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 463:21]
  wire [27:0] ConfigMem_io_out_0; // @[Interconnect.scala 463:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_6_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_7_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_10_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_11_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_out; // @[Interconnect.scala 473:25]
  wire  _T_1 = 10'h5c == io_cfg_addr[11:2]; // @[Interconnect.scala 464:50]
  reg [31:0] _T_12; // @[Interconnect.scala 477:55]
  reg [31:0] _T_14; // @[Interconnect.scala 477:55]
  reg [31:0] _T_16; // @[Interconnect.scala 477:55]
  reg [31:0] _T_18; // @[Interconnect.scala 477:55]
  ConfigMem_90 ConfigMem ( // @[Interconnect.scala 463:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_148 Muxn ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_out(Muxn_io_out)
  );
  Muxn_148 Muxn_1 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_out(Muxn_1_io_out)
  );
  Muxn_148 Muxn_2 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_in_3(Muxn_2_io_in_3),
    .io_out(Muxn_2_io_out)
  );
  Muxn_148 Muxn_3 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_in_3(Muxn_3_io_in_3),
    .io_out(Muxn_3_io_out)
  );
  Muxn_148 Muxn_4 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_in_3(Muxn_4_io_in_3),
    .io_out(Muxn_4_io_out)
  );
  Muxn_148 Muxn_5 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_in_3(Muxn_5_io_in_3),
    .io_out(Muxn_5_io_out)
  );
  Muxn_148 Muxn_6 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_out(Muxn_6_io_out)
  );
  Muxn_148 Muxn_7 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_out(Muxn_7_io_out)
  );
  Muxn_147 Muxn_8 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_147 Muxn_9 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  Muxn_147 Muxn_10 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_10_io_config),
    .io_in_0(Muxn_10_io_in_0),
    .io_in_1(Muxn_10_io_in_1),
    .io_in_2(Muxn_10_io_in_2),
    .io_in_3(Muxn_10_io_in_3),
    .io_in_4(Muxn_10_io_in_4),
    .io_out(Muxn_10_io_out)
  );
  Muxn_147 Muxn_11 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_11_io_config),
    .io_in_0(Muxn_11_io_in_0),
    .io_in_1(Muxn_11_io_in_1),
    .io_in_2(Muxn_11_io_in_2),
    .io_in_3(Muxn_11_io_in_3),
    .io_in_4(Muxn_11_io_in_4),
    .io_out(Muxn_11_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNE_0 = Muxn_2_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinNE_1 = Muxn_3_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinSE_0 = Muxn_4_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSE_1 = Muxn_5_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSW_0 = Muxn_6_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_ipinSW_1 = Muxn_7_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_otrackW_0 = _T_12; // @[Interconnect.scala 430:21 Interconnect.scala 477:45]
  assign io_otrackN_0 = _T_14; // @[Interconnect.scala 431:21 Interconnect.scala 477:45]
  assign io_otrackE_0 = _T_16; // @[Interconnect.scala 432:21 Interconnect.scala 477:45]
  assign io_otrackS_0 = _T_18; // @[Interconnect.scala 433:21 Interconnect.scala 477:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 464:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 466:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 483:23]
  assign Muxn_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 483:23]
  assign Muxn_1_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 483:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 483:23]
  assign Muxn_3_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 483:23]
  assign Muxn_4_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 483:23]
  assign Muxn_5_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[13:12]; // @[Interconnect.scala 483:23]
  assign Muxn_6_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[15:14]; // @[Interconnect.scala 483:23]
  assign Muxn_7_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[18:16]; // @[Interconnect.scala 483:23]
  assign Muxn_8_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[21:19]; // @[Interconnect.scala 483:23]
  assign Muxn_9_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_config = ConfigMem_io_out_0[24:22]; // @[Interconnect.scala 483:23]
  assign Muxn_10_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_config = ConfigMem_io_out_0[27:25]; // @[Interconnect.scala 483:23]
  assign Muxn_11_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_4 = io_itrackE_0; // @[Interconnect.scala 475:63]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_12 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  _T_14 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  _T_16 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  _T_18 = _RAND_3[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_12 <= Muxn_8_io_out;
    _T_14 <= Muxn_9_io_out;
    _T_16 <= Muxn_10_io_out;
    _T_18 <= Muxn_11_io_out;
  end
endmodule
module GIB_38(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
  wire  ConfigMem_clock; // @[Interconnect.scala 463:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 463:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 463:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 463:21]
  wire [27:0] ConfigMem_io_out_0; // @[Interconnect.scala 463:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_6_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_7_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_10_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_11_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_out; // @[Interconnect.scala 473:25]
  wire  _T_1 = 10'h5d == io_cfg_addr[11:2]; // @[Interconnect.scala 464:50]
  ConfigMem_90 ConfigMem ( // @[Interconnect.scala 463:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_148 Muxn ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_out(Muxn_io_out)
  );
  Muxn_148 Muxn_1 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_out(Muxn_1_io_out)
  );
  Muxn_148 Muxn_2 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_in_3(Muxn_2_io_in_3),
    .io_out(Muxn_2_io_out)
  );
  Muxn_148 Muxn_3 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_in_3(Muxn_3_io_in_3),
    .io_out(Muxn_3_io_out)
  );
  Muxn_148 Muxn_4 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_in_3(Muxn_4_io_in_3),
    .io_out(Muxn_4_io_out)
  );
  Muxn_148 Muxn_5 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_in_3(Muxn_5_io_in_3),
    .io_out(Muxn_5_io_out)
  );
  Muxn_148 Muxn_6 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_out(Muxn_6_io_out)
  );
  Muxn_148 Muxn_7 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_out(Muxn_7_io_out)
  );
  Muxn_147 Muxn_8 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_147 Muxn_9 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  Muxn_147 Muxn_10 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_10_io_config),
    .io_in_0(Muxn_10_io_in_0),
    .io_in_1(Muxn_10_io_in_1),
    .io_in_2(Muxn_10_io_in_2),
    .io_in_3(Muxn_10_io_in_3),
    .io_in_4(Muxn_10_io_in_4),
    .io_out(Muxn_10_io_out)
  );
  Muxn_147 Muxn_11 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_11_io_config),
    .io_in_0(Muxn_11_io_in_0),
    .io_in_1(Muxn_11_io_in_1),
    .io_in_2(Muxn_11_io_in_2),
    .io_in_3(Muxn_11_io_in_3),
    .io_in_4(Muxn_11_io_in_4),
    .io_out(Muxn_11_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNE_0 = Muxn_2_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinNE_1 = Muxn_3_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinSE_0 = Muxn_4_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSE_1 = Muxn_5_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSW_0 = Muxn_6_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_ipinSW_1 = Muxn_7_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_otrackW_0 = Muxn_8_io_out; // @[Interconnect.scala 430:21 Interconnect.scala 479:45]
  assign io_otrackN_0 = Muxn_9_io_out; // @[Interconnect.scala 431:21 Interconnect.scala 479:45]
  assign io_otrackE_0 = Muxn_10_io_out; // @[Interconnect.scala 432:21 Interconnect.scala 479:45]
  assign io_otrackS_0 = Muxn_11_io_out; // @[Interconnect.scala 433:21 Interconnect.scala 479:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 464:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 466:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 483:23]
  assign Muxn_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 483:23]
  assign Muxn_1_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 483:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 483:23]
  assign Muxn_3_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 483:23]
  assign Muxn_4_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 483:23]
  assign Muxn_5_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[13:12]; // @[Interconnect.scala 483:23]
  assign Muxn_6_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[15:14]; // @[Interconnect.scala 483:23]
  assign Muxn_7_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[18:16]; // @[Interconnect.scala 483:23]
  assign Muxn_8_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[21:19]; // @[Interconnect.scala 483:23]
  assign Muxn_9_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_config = ConfigMem_io_out_0[24:22]; // @[Interconnect.scala 483:23]
  assign Muxn_10_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_config = ConfigMem_io_out_0[27:25]; // @[Interconnect.scala 483:23]
  assign Muxn_11_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_4 = io_itrackE_0; // @[Interconnect.scala 475:63]
endmodule
module GIB_39(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire  ConfigMem_clock; // @[Interconnect.scala 463:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 463:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 463:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 463:21]
  wire [27:0] ConfigMem_io_out_0; // @[Interconnect.scala 463:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_6_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_7_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_10_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_11_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_out; // @[Interconnect.scala 473:25]
  wire  _T_1 = 10'h5e == io_cfg_addr[11:2]; // @[Interconnect.scala 464:50]
  reg [31:0] _T_12; // @[Interconnect.scala 477:55]
  reg [31:0] _T_14; // @[Interconnect.scala 477:55]
  reg [31:0] _T_16; // @[Interconnect.scala 477:55]
  reg [31:0] _T_18; // @[Interconnect.scala 477:55]
  ConfigMem_90 ConfigMem ( // @[Interconnect.scala 463:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_148 Muxn ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_out(Muxn_io_out)
  );
  Muxn_148 Muxn_1 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_out(Muxn_1_io_out)
  );
  Muxn_148 Muxn_2 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_in_3(Muxn_2_io_in_3),
    .io_out(Muxn_2_io_out)
  );
  Muxn_148 Muxn_3 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_in_3(Muxn_3_io_in_3),
    .io_out(Muxn_3_io_out)
  );
  Muxn_148 Muxn_4 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_in_3(Muxn_4_io_in_3),
    .io_out(Muxn_4_io_out)
  );
  Muxn_148 Muxn_5 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_in_3(Muxn_5_io_in_3),
    .io_out(Muxn_5_io_out)
  );
  Muxn_148 Muxn_6 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_out(Muxn_6_io_out)
  );
  Muxn_148 Muxn_7 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_out(Muxn_7_io_out)
  );
  Muxn_147 Muxn_8 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_147 Muxn_9 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  Muxn_147 Muxn_10 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_10_io_config),
    .io_in_0(Muxn_10_io_in_0),
    .io_in_1(Muxn_10_io_in_1),
    .io_in_2(Muxn_10_io_in_2),
    .io_in_3(Muxn_10_io_in_3),
    .io_in_4(Muxn_10_io_in_4),
    .io_out(Muxn_10_io_out)
  );
  Muxn_147 Muxn_11 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_11_io_config),
    .io_in_0(Muxn_11_io_in_0),
    .io_in_1(Muxn_11_io_in_1),
    .io_in_2(Muxn_11_io_in_2),
    .io_in_3(Muxn_11_io_in_3),
    .io_in_4(Muxn_11_io_in_4),
    .io_out(Muxn_11_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNE_0 = Muxn_2_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinNE_1 = Muxn_3_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinSE_0 = Muxn_4_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSE_1 = Muxn_5_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSW_0 = Muxn_6_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_ipinSW_1 = Muxn_7_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_otrackW_0 = _T_12; // @[Interconnect.scala 430:21 Interconnect.scala 477:45]
  assign io_otrackN_0 = _T_14; // @[Interconnect.scala 431:21 Interconnect.scala 477:45]
  assign io_otrackE_0 = _T_16; // @[Interconnect.scala 432:21 Interconnect.scala 477:45]
  assign io_otrackS_0 = _T_18; // @[Interconnect.scala 433:21 Interconnect.scala 477:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 464:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 466:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 483:23]
  assign Muxn_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 483:23]
  assign Muxn_1_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 483:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 483:23]
  assign Muxn_3_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 483:23]
  assign Muxn_4_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 483:23]
  assign Muxn_5_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[13:12]; // @[Interconnect.scala 483:23]
  assign Muxn_6_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[15:14]; // @[Interconnect.scala 483:23]
  assign Muxn_7_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[18:16]; // @[Interconnect.scala 483:23]
  assign Muxn_8_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[21:19]; // @[Interconnect.scala 483:23]
  assign Muxn_9_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_config = ConfigMem_io_out_0[24:22]; // @[Interconnect.scala 483:23]
  assign Muxn_10_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_config = ConfigMem_io_out_0[27:25]; // @[Interconnect.scala 483:23]
  assign Muxn_11_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_4 = io_itrackE_0; // @[Interconnect.scala 475:63]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_12 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  _T_14 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  _T_16 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  _T_18 = _RAND_3[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_12 <= Muxn_8_io_out;
    _T_14 <= Muxn_9_io_out;
    _T_16 <= Muxn_10_io_out;
    _T_18 <= Muxn_11_io_out;
  end
endmodule
module GIB_40(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
  wire  ConfigMem_clock; // @[Interconnect.scala 463:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 463:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 463:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 463:21]
  wire [27:0] ConfigMem_io_out_0; // @[Interconnect.scala 463:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_6_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_7_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_10_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_11_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_out; // @[Interconnect.scala 473:25]
  wire  _T_1 = 10'h5f == io_cfg_addr[11:2]; // @[Interconnect.scala 464:50]
  ConfigMem_90 ConfigMem ( // @[Interconnect.scala 463:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_148 Muxn ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_out(Muxn_io_out)
  );
  Muxn_148 Muxn_1 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_out(Muxn_1_io_out)
  );
  Muxn_148 Muxn_2 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_in_3(Muxn_2_io_in_3),
    .io_out(Muxn_2_io_out)
  );
  Muxn_148 Muxn_3 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_in_3(Muxn_3_io_in_3),
    .io_out(Muxn_3_io_out)
  );
  Muxn_148 Muxn_4 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_in_3(Muxn_4_io_in_3),
    .io_out(Muxn_4_io_out)
  );
  Muxn_148 Muxn_5 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_in_3(Muxn_5_io_in_3),
    .io_out(Muxn_5_io_out)
  );
  Muxn_148 Muxn_6 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_out(Muxn_6_io_out)
  );
  Muxn_148 Muxn_7 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_out(Muxn_7_io_out)
  );
  Muxn_147 Muxn_8 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_147 Muxn_9 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  Muxn_147 Muxn_10 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_10_io_config),
    .io_in_0(Muxn_10_io_in_0),
    .io_in_1(Muxn_10_io_in_1),
    .io_in_2(Muxn_10_io_in_2),
    .io_in_3(Muxn_10_io_in_3),
    .io_in_4(Muxn_10_io_in_4),
    .io_out(Muxn_10_io_out)
  );
  Muxn_147 Muxn_11 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_11_io_config),
    .io_in_0(Muxn_11_io_in_0),
    .io_in_1(Muxn_11_io_in_1),
    .io_in_2(Muxn_11_io_in_2),
    .io_in_3(Muxn_11_io_in_3),
    .io_in_4(Muxn_11_io_in_4),
    .io_out(Muxn_11_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNE_0 = Muxn_2_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinNE_1 = Muxn_3_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinSE_0 = Muxn_4_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSE_1 = Muxn_5_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSW_0 = Muxn_6_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_ipinSW_1 = Muxn_7_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_otrackW_0 = Muxn_8_io_out; // @[Interconnect.scala 430:21 Interconnect.scala 479:45]
  assign io_otrackN_0 = Muxn_9_io_out; // @[Interconnect.scala 431:21 Interconnect.scala 479:45]
  assign io_otrackE_0 = Muxn_10_io_out; // @[Interconnect.scala 432:21 Interconnect.scala 479:45]
  assign io_otrackS_0 = Muxn_11_io_out; // @[Interconnect.scala 433:21 Interconnect.scala 479:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 464:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 466:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 483:23]
  assign Muxn_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 483:23]
  assign Muxn_1_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 483:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 483:23]
  assign Muxn_3_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 483:23]
  assign Muxn_4_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 483:23]
  assign Muxn_5_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[13:12]; // @[Interconnect.scala 483:23]
  assign Muxn_6_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[15:14]; // @[Interconnect.scala 483:23]
  assign Muxn_7_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[18:16]; // @[Interconnect.scala 483:23]
  assign Muxn_8_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[21:19]; // @[Interconnect.scala 483:23]
  assign Muxn_9_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_config = ConfigMem_io_out_0[24:22]; // @[Interconnect.scala 483:23]
  assign Muxn_10_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_config = ConfigMem_io_out_0[27:25]; // @[Interconnect.scala 483:23]
  assign Muxn_11_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_4 = io_itrackE_0; // @[Interconnect.scala 475:63]
endmodule
module GIB_41(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire  ConfigMem_clock; // @[Interconnect.scala 463:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 463:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 463:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 463:21]
  wire [27:0] ConfigMem_io_out_0; // @[Interconnect.scala 463:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_6_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_7_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_10_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_11_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_out; // @[Interconnect.scala 473:25]
  wire  _T_1 = 10'h60 == io_cfg_addr[11:2]; // @[Interconnect.scala 464:50]
  reg [31:0] _T_12; // @[Interconnect.scala 477:55]
  reg [31:0] _T_14; // @[Interconnect.scala 477:55]
  reg [31:0] _T_16; // @[Interconnect.scala 477:55]
  reg [31:0] _T_18; // @[Interconnect.scala 477:55]
  ConfigMem_90 ConfigMem ( // @[Interconnect.scala 463:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_148 Muxn ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_out(Muxn_io_out)
  );
  Muxn_148 Muxn_1 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_out(Muxn_1_io_out)
  );
  Muxn_148 Muxn_2 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_in_3(Muxn_2_io_in_3),
    .io_out(Muxn_2_io_out)
  );
  Muxn_148 Muxn_3 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_in_3(Muxn_3_io_in_3),
    .io_out(Muxn_3_io_out)
  );
  Muxn_148 Muxn_4 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_in_3(Muxn_4_io_in_3),
    .io_out(Muxn_4_io_out)
  );
  Muxn_148 Muxn_5 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_in_3(Muxn_5_io_in_3),
    .io_out(Muxn_5_io_out)
  );
  Muxn_148 Muxn_6 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_out(Muxn_6_io_out)
  );
  Muxn_148 Muxn_7 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_out(Muxn_7_io_out)
  );
  Muxn_147 Muxn_8 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_147 Muxn_9 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  Muxn_147 Muxn_10 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_10_io_config),
    .io_in_0(Muxn_10_io_in_0),
    .io_in_1(Muxn_10_io_in_1),
    .io_in_2(Muxn_10_io_in_2),
    .io_in_3(Muxn_10_io_in_3),
    .io_in_4(Muxn_10_io_in_4),
    .io_out(Muxn_10_io_out)
  );
  Muxn_147 Muxn_11 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_11_io_config),
    .io_in_0(Muxn_11_io_in_0),
    .io_in_1(Muxn_11_io_in_1),
    .io_in_2(Muxn_11_io_in_2),
    .io_in_3(Muxn_11_io_in_3),
    .io_in_4(Muxn_11_io_in_4),
    .io_out(Muxn_11_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNE_0 = Muxn_2_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinNE_1 = Muxn_3_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinSE_0 = Muxn_4_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSE_1 = Muxn_5_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSW_0 = Muxn_6_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_ipinSW_1 = Muxn_7_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_otrackW_0 = _T_12; // @[Interconnect.scala 430:21 Interconnect.scala 477:45]
  assign io_otrackN_0 = _T_14; // @[Interconnect.scala 431:21 Interconnect.scala 477:45]
  assign io_otrackE_0 = _T_16; // @[Interconnect.scala 432:21 Interconnect.scala 477:45]
  assign io_otrackS_0 = _T_18; // @[Interconnect.scala 433:21 Interconnect.scala 477:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 464:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 466:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 483:23]
  assign Muxn_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 483:23]
  assign Muxn_1_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 483:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 483:23]
  assign Muxn_3_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 483:23]
  assign Muxn_4_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 483:23]
  assign Muxn_5_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[13:12]; // @[Interconnect.scala 483:23]
  assign Muxn_6_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[15:14]; // @[Interconnect.scala 483:23]
  assign Muxn_7_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[18:16]; // @[Interconnect.scala 483:23]
  assign Muxn_8_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[21:19]; // @[Interconnect.scala 483:23]
  assign Muxn_9_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_config = ConfigMem_io_out_0[24:22]; // @[Interconnect.scala 483:23]
  assign Muxn_10_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_config = ConfigMem_io_out_0[27:25]; // @[Interconnect.scala 483:23]
  assign Muxn_11_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_4 = io_itrackE_0; // @[Interconnect.scala 475:63]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_12 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  _T_14 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  _T_16 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  _T_18 = _RAND_3[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_12 <= Muxn_8_io_out;
    _T_14 <= Muxn_9_io_out;
    _T_16 <= Muxn_10_io_out;
    _T_18 <= Muxn_11_io_out;
  end
endmodule
module GIB_42(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
  wire  ConfigMem_clock; // @[Interconnect.scala 463:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 463:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 463:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 463:21]
  wire [27:0] ConfigMem_io_out_0; // @[Interconnect.scala 463:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_6_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_7_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_10_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_11_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_out; // @[Interconnect.scala 473:25]
  wire  _T_1 = 10'h61 == io_cfg_addr[11:2]; // @[Interconnect.scala 464:50]
  ConfigMem_90 ConfigMem ( // @[Interconnect.scala 463:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_148 Muxn ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_out(Muxn_io_out)
  );
  Muxn_148 Muxn_1 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_out(Muxn_1_io_out)
  );
  Muxn_148 Muxn_2 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_in_3(Muxn_2_io_in_3),
    .io_out(Muxn_2_io_out)
  );
  Muxn_148 Muxn_3 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_in_3(Muxn_3_io_in_3),
    .io_out(Muxn_3_io_out)
  );
  Muxn_148 Muxn_4 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_in_3(Muxn_4_io_in_3),
    .io_out(Muxn_4_io_out)
  );
  Muxn_148 Muxn_5 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_in_3(Muxn_5_io_in_3),
    .io_out(Muxn_5_io_out)
  );
  Muxn_148 Muxn_6 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_out(Muxn_6_io_out)
  );
  Muxn_148 Muxn_7 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_out(Muxn_7_io_out)
  );
  Muxn_147 Muxn_8 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_147 Muxn_9 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  Muxn_147 Muxn_10 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_10_io_config),
    .io_in_0(Muxn_10_io_in_0),
    .io_in_1(Muxn_10_io_in_1),
    .io_in_2(Muxn_10_io_in_2),
    .io_in_3(Muxn_10_io_in_3),
    .io_in_4(Muxn_10_io_in_4),
    .io_out(Muxn_10_io_out)
  );
  Muxn_147 Muxn_11 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_11_io_config),
    .io_in_0(Muxn_11_io_in_0),
    .io_in_1(Muxn_11_io_in_1),
    .io_in_2(Muxn_11_io_in_2),
    .io_in_3(Muxn_11_io_in_3),
    .io_in_4(Muxn_11_io_in_4),
    .io_out(Muxn_11_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNE_0 = Muxn_2_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinNE_1 = Muxn_3_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinSE_0 = Muxn_4_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSE_1 = Muxn_5_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSW_0 = Muxn_6_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_ipinSW_1 = Muxn_7_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_otrackW_0 = Muxn_8_io_out; // @[Interconnect.scala 430:21 Interconnect.scala 479:45]
  assign io_otrackN_0 = Muxn_9_io_out; // @[Interconnect.scala 431:21 Interconnect.scala 479:45]
  assign io_otrackE_0 = Muxn_10_io_out; // @[Interconnect.scala 432:21 Interconnect.scala 479:45]
  assign io_otrackS_0 = Muxn_11_io_out; // @[Interconnect.scala 433:21 Interconnect.scala 479:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 464:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 466:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 483:23]
  assign Muxn_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 483:23]
  assign Muxn_1_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 483:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 483:23]
  assign Muxn_3_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 483:23]
  assign Muxn_4_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 483:23]
  assign Muxn_5_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[13:12]; // @[Interconnect.scala 483:23]
  assign Muxn_6_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[15:14]; // @[Interconnect.scala 483:23]
  assign Muxn_7_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[18:16]; // @[Interconnect.scala 483:23]
  assign Muxn_8_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[21:19]; // @[Interconnect.scala 483:23]
  assign Muxn_9_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_config = ConfigMem_io_out_0[24:22]; // @[Interconnect.scala 483:23]
  assign Muxn_10_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_config = ConfigMem_io_out_0[27:25]; // @[Interconnect.scala 483:23]
  assign Muxn_11_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_4 = io_itrackE_0; // @[Interconnect.scala 475:63]
endmodule
module GIB_43(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire  ConfigMem_clock; // @[Interconnect.scala 463:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 463:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 463:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 463:21]
  wire [27:0] ConfigMem_io_out_0; // @[Interconnect.scala 463:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_6_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_7_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_10_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_11_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_out; // @[Interconnect.scala 473:25]
  wire  _T_1 = 10'h62 == io_cfg_addr[11:2]; // @[Interconnect.scala 464:50]
  reg [31:0] _T_12; // @[Interconnect.scala 477:55]
  reg [31:0] _T_14; // @[Interconnect.scala 477:55]
  reg [31:0] _T_16; // @[Interconnect.scala 477:55]
  reg [31:0] _T_18; // @[Interconnect.scala 477:55]
  ConfigMem_90 ConfigMem ( // @[Interconnect.scala 463:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_148 Muxn ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_out(Muxn_io_out)
  );
  Muxn_148 Muxn_1 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_out(Muxn_1_io_out)
  );
  Muxn_148 Muxn_2 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_in_3(Muxn_2_io_in_3),
    .io_out(Muxn_2_io_out)
  );
  Muxn_148 Muxn_3 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_in_3(Muxn_3_io_in_3),
    .io_out(Muxn_3_io_out)
  );
  Muxn_148 Muxn_4 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_in_3(Muxn_4_io_in_3),
    .io_out(Muxn_4_io_out)
  );
  Muxn_148 Muxn_5 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_in_3(Muxn_5_io_in_3),
    .io_out(Muxn_5_io_out)
  );
  Muxn_148 Muxn_6 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_out(Muxn_6_io_out)
  );
  Muxn_148 Muxn_7 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_out(Muxn_7_io_out)
  );
  Muxn_147 Muxn_8 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_147 Muxn_9 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  Muxn_147 Muxn_10 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_10_io_config),
    .io_in_0(Muxn_10_io_in_0),
    .io_in_1(Muxn_10_io_in_1),
    .io_in_2(Muxn_10_io_in_2),
    .io_in_3(Muxn_10_io_in_3),
    .io_in_4(Muxn_10_io_in_4),
    .io_out(Muxn_10_io_out)
  );
  Muxn_147 Muxn_11 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_11_io_config),
    .io_in_0(Muxn_11_io_in_0),
    .io_in_1(Muxn_11_io_in_1),
    .io_in_2(Muxn_11_io_in_2),
    .io_in_3(Muxn_11_io_in_3),
    .io_in_4(Muxn_11_io_in_4),
    .io_out(Muxn_11_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNE_0 = Muxn_2_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinNE_1 = Muxn_3_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinSE_0 = Muxn_4_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSE_1 = Muxn_5_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSW_0 = Muxn_6_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_ipinSW_1 = Muxn_7_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_otrackW_0 = _T_12; // @[Interconnect.scala 430:21 Interconnect.scala 477:45]
  assign io_otrackN_0 = _T_14; // @[Interconnect.scala 431:21 Interconnect.scala 477:45]
  assign io_otrackE_0 = _T_16; // @[Interconnect.scala 432:21 Interconnect.scala 477:45]
  assign io_otrackS_0 = _T_18; // @[Interconnect.scala 433:21 Interconnect.scala 477:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 464:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 466:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 483:23]
  assign Muxn_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 483:23]
  assign Muxn_1_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 483:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 483:23]
  assign Muxn_3_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 483:23]
  assign Muxn_4_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 483:23]
  assign Muxn_5_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[13:12]; // @[Interconnect.scala 483:23]
  assign Muxn_6_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[15:14]; // @[Interconnect.scala 483:23]
  assign Muxn_7_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[18:16]; // @[Interconnect.scala 483:23]
  assign Muxn_8_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[21:19]; // @[Interconnect.scala 483:23]
  assign Muxn_9_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_config = ConfigMem_io_out_0[24:22]; // @[Interconnect.scala 483:23]
  assign Muxn_10_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_config = ConfigMem_io_out_0[27:25]; // @[Interconnect.scala 483:23]
  assign Muxn_11_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_4 = io_itrackE_0; // @[Interconnect.scala 475:63]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_12 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  _T_14 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  _T_16 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  _T_18 = _RAND_3[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_12 <= Muxn_8_io_out;
    _T_14 <= Muxn_9_io_out;
    _T_16 <= Muxn_10_io_out;
    _T_18 <= Muxn_11_io_out;
  end
endmodule
module GIB_44(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
  wire  ConfigMem_clock; // @[Interconnect.scala 463:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 463:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 463:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 463:21]
  wire [14:0] ConfigMem_io_out_0; // @[Interconnect.scala 463:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 473:25]
  wire  Muxn_2_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 473:25]
  wire  Muxn_3_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_6_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_7_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 473:25]
  wire  _T_1 = 10'h63 == io_cfg_addr[11:2]; // @[Interconnect.scala 464:50]
  ConfigMem_89 ConfigMem ( // @[Interconnect.scala 463:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_145 Muxn ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_out(Muxn_io_out)
  );
  Muxn_145 Muxn_1 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_out(Muxn_1_io_out)
  );
  Muxn Muxn_2 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_out(Muxn_2_io_out)
  );
  Muxn Muxn_3 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_out(Muxn_3_io_out)
  );
  Muxn_145 Muxn_4 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_out(Muxn_4_io_out)
  );
  Muxn_148 Muxn_5 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_in_3(Muxn_5_io_in_3),
    .io_out(Muxn_5_io_out)
  );
  Muxn_147 Muxn_6 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_in_4(Muxn_6_io_in_4),
    .io_out(Muxn_6_io_out)
  );
  Muxn_148 Muxn_7 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_out(Muxn_7_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinSW_0 = Muxn_2_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_ipinSW_1 = Muxn_3_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_otrackW_0 = Muxn_4_io_out; // @[Interconnect.scala 430:21 Interconnect.scala 479:45]
  assign io_otrackN_0 = Muxn_5_io_out; // @[Interconnect.scala 431:21 Interconnect.scala 479:45]
  assign io_otrackS_0 = Muxn_7_io_out; // @[Interconnect.scala 433:21 Interconnect.scala 479:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 464:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 466:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 483:23]
  assign Muxn_io_in_0 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_1 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_2 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 483:23]
  assign Muxn_1_io_in_0 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_1 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_2 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[4]; // @[Interconnect.scala 483:23]
  assign Muxn_2_io_in_0 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_1 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[5]; // @[Interconnect.scala 483:23]
  assign Muxn_3_io_in_0 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_1 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 483:23]
  assign Muxn_4_io_in_0 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_1 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_2 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 483:23]
  assign Muxn_5_io_in_0 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_1 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_2 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[12:10]; // @[Interconnect.scala 483:23]
  assign Muxn_6_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[14:13]; // @[Interconnect.scala 483:23]
  assign Muxn_7_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_1 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_3 = 32'h0; // @[Interconnect.scala 475:63]
endmodule
module GIB_45(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire  ConfigMem_clock; // @[Interconnect.scala 463:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 463:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 463:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 463:21]
  wire [14:0] ConfigMem_io_out_0; // @[Interconnect.scala 463:21]
  wire  Muxn_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 473:25]
  wire  Muxn_1_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_4_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_6_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_7_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 473:25]
  wire  _T_1 = 10'h6d == io_cfg_addr[11:2]; // @[Interconnect.scala 464:50]
  reg [31:0] _T_10; // @[Interconnect.scala 477:55]
  reg [31:0] _T_12; // @[Interconnect.scala 477:55]
  reg [31:0] _T_14; // @[Interconnect.scala 477:55]
  ConfigMem_89 ConfigMem ( // @[Interconnect.scala 463:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn Muxn ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_out(Muxn_io_out)
  );
  Muxn Muxn_1 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_out(Muxn_1_io_out)
  );
  Muxn_145 Muxn_2 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_out(Muxn_2_io_out)
  );
  Muxn_145 Muxn_3 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_out(Muxn_3_io_out)
  );
  Muxn_147 Muxn_4 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_in_3(Muxn_4_io_in_3),
    .io_in_4(Muxn_4_io_in_4),
    .io_out(Muxn_4_io_out)
  );
  Muxn_148 Muxn_5 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_in_3(Muxn_5_io_in_3),
    .io_out(Muxn_5_io_out)
  );
  Muxn_145 Muxn_6 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_out(Muxn_6_io_out)
  );
  Muxn_148 Muxn_7 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_out(Muxn_7_io_out)
  );
  assign io_ipinNE_0 = Muxn_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinNE_1 = Muxn_1_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinSE_0 = Muxn_2_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSE_1 = Muxn_3_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_otrackN_0 = _T_10; // @[Interconnect.scala 431:21 Interconnect.scala 477:45]
  assign io_otrackE_0 = _T_12; // @[Interconnect.scala 432:21 Interconnect.scala 477:45]
  assign io_otrackS_0 = _T_14; // @[Interconnect.scala 433:21 Interconnect.scala 477:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 464:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 466:21]
  assign Muxn_io_config = ConfigMem_io_out_0[0]; // @[Interconnect.scala 483:23]
  assign Muxn_io_in_0 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_1 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[1]; // @[Interconnect.scala 483:23]
  assign Muxn_1_io_in_0 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_1 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 483:23]
  assign Muxn_2_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_1 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 483:23]
  assign Muxn_3_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_1 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[8:6]; // @[Interconnect.scala 483:23]
  assign Muxn_4_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[10:9]; // @[Interconnect.scala 483:23]
  assign Muxn_5_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_1 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[12:11]; // @[Interconnect.scala 483:23]
  assign Muxn_6_io_in_0 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_1 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_2 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[14:13]; // @[Interconnect.scala 483:23]
  assign Muxn_7_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_1 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_10 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  _T_12 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  _T_14 = _RAND_2[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_10 <= Muxn_5_io_out;
    _T_12 <= Muxn_6_io_out;
    _T_14 <= Muxn_7_io_out;
  end
endmodule
module GIB_46(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
  wire  ConfigMem_clock; // @[Interconnect.scala 463:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 463:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 463:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 463:21]
  wire [27:0] ConfigMem_io_out_0; // @[Interconnect.scala 463:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_6_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_7_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_10_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_11_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_out; // @[Interconnect.scala 473:25]
  wire  _T_1 = 10'h6e == io_cfg_addr[11:2]; // @[Interconnect.scala 464:50]
  ConfigMem_90 ConfigMem ( // @[Interconnect.scala 463:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_148 Muxn ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_out(Muxn_io_out)
  );
  Muxn_148 Muxn_1 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_out(Muxn_1_io_out)
  );
  Muxn_148 Muxn_2 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_in_3(Muxn_2_io_in_3),
    .io_out(Muxn_2_io_out)
  );
  Muxn_148 Muxn_3 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_in_3(Muxn_3_io_in_3),
    .io_out(Muxn_3_io_out)
  );
  Muxn_148 Muxn_4 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_in_3(Muxn_4_io_in_3),
    .io_out(Muxn_4_io_out)
  );
  Muxn_148 Muxn_5 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_in_3(Muxn_5_io_in_3),
    .io_out(Muxn_5_io_out)
  );
  Muxn_148 Muxn_6 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_out(Muxn_6_io_out)
  );
  Muxn_148 Muxn_7 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_out(Muxn_7_io_out)
  );
  Muxn_147 Muxn_8 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_147 Muxn_9 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  Muxn_147 Muxn_10 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_10_io_config),
    .io_in_0(Muxn_10_io_in_0),
    .io_in_1(Muxn_10_io_in_1),
    .io_in_2(Muxn_10_io_in_2),
    .io_in_3(Muxn_10_io_in_3),
    .io_in_4(Muxn_10_io_in_4),
    .io_out(Muxn_10_io_out)
  );
  Muxn_147 Muxn_11 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_11_io_config),
    .io_in_0(Muxn_11_io_in_0),
    .io_in_1(Muxn_11_io_in_1),
    .io_in_2(Muxn_11_io_in_2),
    .io_in_3(Muxn_11_io_in_3),
    .io_in_4(Muxn_11_io_in_4),
    .io_out(Muxn_11_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNE_0 = Muxn_2_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinNE_1 = Muxn_3_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinSE_0 = Muxn_4_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSE_1 = Muxn_5_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSW_0 = Muxn_6_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_ipinSW_1 = Muxn_7_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_otrackW_0 = Muxn_8_io_out; // @[Interconnect.scala 430:21 Interconnect.scala 479:45]
  assign io_otrackN_0 = Muxn_9_io_out; // @[Interconnect.scala 431:21 Interconnect.scala 479:45]
  assign io_otrackE_0 = Muxn_10_io_out; // @[Interconnect.scala 432:21 Interconnect.scala 479:45]
  assign io_otrackS_0 = Muxn_11_io_out; // @[Interconnect.scala 433:21 Interconnect.scala 479:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 464:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 466:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 483:23]
  assign Muxn_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 483:23]
  assign Muxn_1_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 483:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 483:23]
  assign Muxn_3_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 483:23]
  assign Muxn_4_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 483:23]
  assign Muxn_5_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[13:12]; // @[Interconnect.scala 483:23]
  assign Muxn_6_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[15:14]; // @[Interconnect.scala 483:23]
  assign Muxn_7_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[18:16]; // @[Interconnect.scala 483:23]
  assign Muxn_8_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[21:19]; // @[Interconnect.scala 483:23]
  assign Muxn_9_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_config = ConfigMem_io_out_0[24:22]; // @[Interconnect.scala 483:23]
  assign Muxn_10_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_config = ConfigMem_io_out_0[27:25]; // @[Interconnect.scala 483:23]
  assign Muxn_11_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_4 = io_itrackE_0; // @[Interconnect.scala 475:63]
endmodule
module GIB_47(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire  ConfigMem_clock; // @[Interconnect.scala 463:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 463:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 463:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 463:21]
  wire [27:0] ConfigMem_io_out_0; // @[Interconnect.scala 463:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_6_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_7_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_10_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_11_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_out; // @[Interconnect.scala 473:25]
  wire  _T_1 = 10'h6f == io_cfg_addr[11:2]; // @[Interconnect.scala 464:50]
  reg [31:0] _T_12; // @[Interconnect.scala 477:55]
  reg [31:0] _T_14; // @[Interconnect.scala 477:55]
  reg [31:0] _T_16; // @[Interconnect.scala 477:55]
  reg [31:0] _T_18; // @[Interconnect.scala 477:55]
  ConfigMem_90 ConfigMem ( // @[Interconnect.scala 463:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_148 Muxn ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_out(Muxn_io_out)
  );
  Muxn_148 Muxn_1 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_out(Muxn_1_io_out)
  );
  Muxn_148 Muxn_2 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_in_3(Muxn_2_io_in_3),
    .io_out(Muxn_2_io_out)
  );
  Muxn_148 Muxn_3 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_in_3(Muxn_3_io_in_3),
    .io_out(Muxn_3_io_out)
  );
  Muxn_148 Muxn_4 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_in_3(Muxn_4_io_in_3),
    .io_out(Muxn_4_io_out)
  );
  Muxn_148 Muxn_5 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_in_3(Muxn_5_io_in_3),
    .io_out(Muxn_5_io_out)
  );
  Muxn_148 Muxn_6 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_out(Muxn_6_io_out)
  );
  Muxn_148 Muxn_7 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_out(Muxn_7_io_out)
  );
  Muxn_147 Muxn_8 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_147 Muxn_9 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  Muxn_147 Muxn_10 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_10_io_config),
    .io_in_0(Muxn_10_io_in_0),
    .io_in_1(Muxn_10_io_in_1),
    .io_in_2(Muxn_10_io_in_2),
    .io_in_3(Muxn_10_io_in_3),
    .io_in_4(Muxn_10_io_in_4),
    .io_out(Muxn_10_io_out)
  );
  Muxn_147 Muxn_11 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_11_io_config),
    .io_in_0(Muxn_11_io_in_0),
    .io_in_1(Muxn_11_io_in_1),
    .io_in_2(Muxn_11_io_in_2),
    .io_in_3(Muxn_11_io_in_3),
    .io_in_4(Muxn_11_io_in_4),
    .io_out(Muxn_11_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNE_0 = Muxn_2_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinNE_1 = Muxn_3_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinSE_0 = Muxn_4_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSE_1 = Muxn_5_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSW_0 = Muxn_6_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_ipinSW_1 = Muxn_7_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_otrackW_0 = _T_12; // @[Interconnect.scala 430:21 Interconnect.scala 477:45]
  assign io_otrackN_0 = _T_14; // @[Interconnect.scala 431:21 Interconnect.scala 477:45]
  assign io_otrackE_0 = _T_16; // @[Interconnect.scala 432:21 Interconnect.scala 477:45]
  assign io_otrackS_0 = _T_18; // @[Interconnect.scala 433:21 Interconnect.scala 477:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 464:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 466:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 483:23]
  assign Muxn_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 483:23]
  assign Muxn_1_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 483:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 483:23]
  assign Muxn_3_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 483:23]
  assign Muxn_4_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 483:23]
  assign Muxn_5_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[13:12]; // @[Interconnect.scala 483:23]
  assign Muxn_6_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[15:14]; // @[Interconnect.scala 483:23]
  assign Muxn_7_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[18:16]; // @[Interconnect.scala 483:23]
  assign Muxn_8_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[21:19]; // @[Interconnect.scala 483:23]
  assign Muxn_9_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_config = ConfigMem_io_out_0[24:22]; // @[Interconnect.scala 483:23]
  assign Muxn_10_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_config = ConfigMem_io_out_0[27:25]; // @[Interconnect.scala 483:23]
  assign Muxn_11_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_4 = io_itrackE_0; // @[Interconnect.scala 475:63]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_12 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  _T_14 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  _T_16 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  _T_18 = _RAND_3[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_12 <= Muxn_8_io_out;
    _T_14 <= Muxn_9_io_out;
    _T_16 <= Muxn_10_io_out;
    _T_18 <= Muxn_11_io_out;
  end
endmodule
module GIB_48(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
  wire  ConfigMem_clock; // @[Interconnect.scala 463:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 463:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 463:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 463:21]
  wire [27:0] ConfigMem_io_out_0; // @[Interconnect.scala 463:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_6_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_7_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_10_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_11_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_out; // @[Interconnect.scala 473:25]
  wire  _T_1 = 10'h70 == io_cfg_addr[11:2]; // @[Interconnect.scala 464:50]
  ConfigMem_90 ConfigMem ( // @[Interconnect.scala 463:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_148 Muxn ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_out(Muxn_io_out)
  );
  Muxn_148 Muxn_1 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_out(Muxn_1_io_out)
  );
  Muxn_148 Muxn_2 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_in_3(Muxn_2_io_in_3),
    .io_out(Muxn_2_io_out)
  );
  Muxn_148 Muxn_3 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_in_3(Muxn_3_io_in_3),
    .io_out(Muxn_3_io_out)
  );
  Muxn_148 Muxn_4 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_in_3(Muxn_4_io_in_3),
    .io_out(Muxn_4_io_out)
  );
  Muxn_148 Muxn_5 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_in_3(Muxn_5_io_in_3),
    .io_out(Muxn_5_io_out)
  );
  Muxn_148 Muxn_6 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_out(Muxn_6_io_out)
  );
  Muxn_148 Muxn_7 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_out(Muxn_7_io_out)
  );
  Muxn_147 Muxn_8 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_147 Muxn_9 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  Muxn_147 Muxn_10 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_10_io_config),
    .io_in_0(Muxn_10_io_in_0),
    .io_in_1(Muxn_10_io_in_1),
    .io_in_2(Muxn_10_io_in_2),
    .io_in_3(Muxn_10_io_in_3),
    .io_in_4(Muxn_10_io_in_4),
    .io_out(Muxn_10_io_out)
  );
  Muxn_147 Muxn_11 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_11_io_config),
    .io_in_0(Muxn_11_io_in_0),
    .io_in_1(Muxn_11_io_in_1),
    .io_in_2(Muxn_11_io_in_2),
    .io_in_3(Muxn_11_io_in_3),
    .io_in_4(Muxn_11_io_in_4),
    .io_out(Muxn_11_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNE_0 = Muxn_2_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinNE_1 = Muxn_3_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinSE_0 = Muxn_4_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSE_1 = Muxn_5_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSW_0 = Muxn_6_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_ipinSW_1 = Muxn_7_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_otrackW_0 = Muxn_8_io_out; // @[Interconnect.scala 430:21 Interconnect.scala 479:45]
  assign io_otrackN_0 = Muxn_9_io_out; // @[Interconnect.scala 431:21 Interconnect.scala 479:45]
  assign io_otrackE_0 = Muxn_10_io_out; // @[Interconnect.scala 432:21 Interconnect.scala 479:45]
  assign io_otrackS_0 = Muxn_11_io_out; // @[Interconnect.scala 433:21 Interconnect.scala 479:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 464:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 466:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 483:23]
  assign Muxn_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 483:23]
  assign Muxn_1_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 483:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 483:23]
  assign Muxn_3_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 483:23]
  assign Muxn_4_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 483:23]
  assign Muxn_5_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[13:12]; // @[Interconnect.scala 483:23]
  assign Muxn_6_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[15:14]; // @[Interconnect.scala 483:23]
  assign Muxn_7_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[18:16]; // @[Interconnect.scala 483:23]
  assign Muxn_8_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[21:19]; // @[Interconnect.scala 483:23]
  assign Muxn_9_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_config = ConfigMem_io_out_0[24:22]; // @[Interconnect.scala 483:23]
  assign Muxn_10_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_config = ConfigMem_io_out_0[27:25]; // @[Interconnect.scala 483:23]
  assign Muxn_11_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_4 = io_itrackE_0; // @[Interconnect.scala 475:63]
endmodule
module GIB_49(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire  ConfigMem_clock; // @[Interconnect.scala 463:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 463:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 463:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 463:21]
  wire [27:0] ConfigMem_io_out_0; // @[Interconnect.scala 463:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_6_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_7_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_10_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_11_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_out; // @[Interconnect.scala 473:25]
  wire  _T_1 = 10'h71 == io_cfg_addr[11:2]; // @[Interconnect.scala 464:50]
  reg [31:0] _T_12; // @[Interconnect.scala 477:55]
  reg [31:0] _T_14; // @[Interconnect.scala 477:55]
  reg [31:0] _T_16; // @[Interconnect.scala 477:55]
  reg [31:0] _T_18; // @[Interconnect.scala 477:55]
  ConfigMem_90 ConfigMem ( // @[Interconnect.scala 463:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_148 Muxn ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_out(Muxn_io_out)
  );
  Muxn_148 Muxn_1 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_out(Muxn_1_io_out)
  );
  Muxn_148 Muxn_2 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_in_3(Muxn_2_io_in_3),
    .io_out(Muxn_2_io_out)
  );
  Muxn_148 Muxn_3 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_in_3(Muxn_3_io_in_3),
    .io_out(Muxn_3_io_out)
  );
  Muxn_148 Muxn_4 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_in_3(Muxn_4_io_in_3),
    .io_out(Muxn_4_io_out)
  );
  Muxn_148 Muxn_5 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_in_3(Muxn_5_io_in_3),
    .io_out(Muxn_5_io_out)
  );
  Muxn_148 Muxn_6 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_out(Muxn_6_io_out)
  );
  Muxn_148 Muxn_7 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_out(Muxn_7_io_out)
  );
  Muxn_147 Muxn_8 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_147 Muxn_9 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  Muxn_147 Muxn_10 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_10_io_config),
    .io_in_0(Muxn_10_io_in_0),
    .io_in_1(Muxn_10_io_in_1),
    .io_in_2(Muxn_10_io_in_2),
    .io_in_3(Muxn_10_io_in_3),
    .io_in_4(Muxn_10_io_in_4),
    .io_out(Muxn_10_io_out)
  );
  Muxn_147 Muxn_11 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_11_io_config),
    .io_in_0(Muxn_11_io_in_0),
    .io_in_1(Muxn_11_io_in_1),
    .io_in_2(Muxn_11_io_in_2),
    .io_in_3(Muxn_11_io_in_3),
    .io_in_4(Muxn_11_io_in_4),
    .io_out(Muxn_11_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNE_0 = Muxn_2_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinNE_1 = Muxn_3_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinSE_0 = Muxn_4_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSE_1 = Muxn_5_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSW_0 = Muxn_6_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_ipinSW_1 = Muxn_7_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_otrackW_0 = _T_12; // @[Interconnect.scala 430:21 Interconnect.scala 477:45]
  assign io_otrackN_0 = _T_14; // @[Interconnect.scala 431:21 Interconnect.scala 477:45]
  assign io_otrackE_0 = _T_16; // @[Interconnect.scala 432:21 Interconnect.scala 477:45]
  assign io_otrackS_0 = _T_18; // @[Interconnect.scala 433:21 Interconnect.scala 477:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 464:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 466:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 483:23]
  assign Muxn_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 483:23]
  assign Muxn_1_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 483:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 483:23]
  assign Muxn_3_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 483:23]
  assign Muxn_4_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 483:23]
  assign Muxn_5_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[13:12]; // @[Interconnect.scala 483:23]
  assign Muxn_6_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[15:14]; // @[Interconnect.scala 483:23]
  assign Muxn_7_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[18:16]; // @[Interconnect.scala 483:23]
  assign Muxn_8_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[21:19]; // @[Interconnect.scala 483:23]
  assign Muxn_9_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_config = ConfigMem_io_out_0[24:22]; // @[Interconnect.scala 483:23]
  assign Muxn_10_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_config = ConfigMem_io_out_0[27:25]; // @[Interconnect.scala 483:23]
  assign Muxn_11_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_4 = io_itrackE_0; // @[Interconnect.scala 475:63]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_12 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  _T_14 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  _T_16 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  _T_18 = _RAND_3[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_12 <= Muxn_8_io_out;
    _T_14 <= Muxn_9_io_out;
    _T_16 <= Muxn_10_io_out;
    _T_18 <= Muxn_11_io_out;
  end
endmodule
module GIB_50(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
  wire  ConfigMem_clock; // @[Interconnect.scala 463:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 463:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 463:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 463:21]
  wire [27:0] ConfigMem_io_out_0; // @[Interconnect.scala 463:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_6_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_7_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_10_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_11_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_out; // @[Interconnect.scala 473:25]
  wire  _T_1 = 10'h72 == io_cfg_addr[11:2]; // @[Interconnect.scala 464:50]
  ConfigMem_90 ConfigMem ( // @[Interconnect.scala 463:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_148 Muxn ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_out(Muxn_io_out)
  );
  Muxn_148 Muxn_1 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_out(Muxn_1_io_out)
  );
  Muxn_148 Muxn_2 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_in_3(Muxn_2_io_in_3),
    .io_out(Muxn_2_io_out)
  );
  Muxn_148 Muxn_3 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_in_3(Muxn_3_io_in_3),
    .io_out(Muxn_3_io_out)
  );
  Muxn_148 Muxn_4 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_in_3(Muxn_4_io_in_3),
    .io_out(Muxn_4_io_out)
  );
  Muxn_148 Muxn_5 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_in_3(Muxn_5_io_in_3),
    .io_out(Muxn_5_io_out)
  );
  Muxn_148 Muxn_6 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_out(Muxn_6_io_out)
  );
  Muxn_148 Muxn_7 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_out(Muxn_7_io_out)
  );
  Muxn_147 Muxn_8 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_147 Muxn_9 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  Muxn_147 Muxn_10 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_10_io_config),
    .io_in_0(Muxn_10_io_in_0),
    .io_in_1(Muxn_10_io_in_1),
    .io_in_2(Muxn_10_io_in_2),
    .io_in_3(Muxn_10_io_in_3),
    .io_in_4(Muxn_10_io_in_4),
    .io_out(Muxn_10_io_out)
  );
  Muxn_147 Muxn_11 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_11_io_config),
    .io_in_0(Muxn_11_io_in_0),
    .io_in_1(Muxn_11_io_in_1),
    .io_in_2(Muxn_11_io_in_2),
    .io_in_3(Muxn_11_io_in_3),
    .io_in_4(Muxn_11_io_in_4),
    .io_out(Muxn_11_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNE_0 = Muxn_2_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinNE_1 = Muxn_3_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinSE_0 = Muxn_4_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSE_1 = Muxn_5_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSW_0 = Muxn_6_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_ipinSW_1 = Muxn_7_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_otrackW_0 = Muxn_8_io_out; // @[Interconnect.scala 430:21 Interconnect.scala 479:45]
  assign io_otrackN_0 = Muxn_9_io_out; // @[Interconnect.scala 431:21 Interconnect.scala 479:45]
  assign io_otrackE_0 = Muxn_10_io_out; // @[Interconnect.scala 432:21 Interconnect.scala 479:45]
  assign io_otrackS_0 = Muxn_11_io_out; // @[Interconnect.scala 433:21 Interconnect.scala 479:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 464:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 466:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 483:23]
  assign Muxn_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 483:23]
  assign Muxn_1_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 483:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 483:23]
  assign Muxn_3_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 483:23]
  assign Muxn_4_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 483:23]
  assign Muxn_5_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[13:12]; // @[Interconnect.scala 483:23]
  assign Muxn_6_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[15:14]; // @[Interconnect.scala 483:23]
  assign Muxn_7_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[18:16]; // @[Interconnect.scala 483:23]
  assign Muxn_8_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[21:19]; // @[Interconnect.scala 483:23]
  assign Muxn_9_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_config = ConfigMem_io_out_0[24:22]; // @[Interconnect.scala 483:23]
  assign Muxn_10_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_config = ConfigMem_io_out_0[27:25]; // @[Interconnect.scala 483:23]
  assign Muxn_11_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_4 = io_itrackE_0; // @[Interconnect.scala 475:63]
endmodule
module GIB_51(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire  ConfigMem_clock; // @[Interconnect.scala 463:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 463:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 463:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 463:21]
  wire [27:0] ConfigMem_io_out_0; // @[Interconnect.scala 463:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_6_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_7_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_10_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_11_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_out; // @[Interconnect.scala 473:25]
  wire  _T_1 = 10'h73 == io_cfg_addr[11:2]; // @[Interconnect.scala 464:50]
  reg [31:0] _T_12; // @[Interconnect.scala 477:55]
  reg [31:0] _T_14; // @[Interconnect.scala 477:55]
  reg [31:0] _T_16; // @[Interconnect.scala 477:55]
  reg [31:0] _T_18; // @[Interconnect.scala 477:55]
  ConfigMem_90 ConfigMem ( // @[Interconnect.scala 463:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_148 Muxn ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_out(Muxn_io_out)
  );
  Muxn_148 Muxn_1 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_out(Muxn_1_io_out)
  );
  Muxn_148 Muxn_2 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_in_3(Muxn_2_io_in_3),
    .io_out(Muxn_2_io_out)
  );
  Muxn_148 Muxn_3 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_in_3(Muxn_3_io_in_3),
    .io_out(Muxn_3_io_out)
  );
  Muxn_148 Muxn_4 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_in_3(Muxn_4_io_in_3),
    .io_out(Muxn_4_io_out)
  );
  Muxn_148 Muxn_5 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_in_3(Muxn_5_io_in_3),
    .io_out(Muxn_5_io_out)
  );
  Muxn_148 Muxn_6 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_out(Muxn_6_io_out)
  );
  Muxn_148 Muxn_7 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_out(Muxn_7_io_out)
  );
  Muxn_147 Muxn_8 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_147 Muxn_9 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  Muxn_147 Muxn_10 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_10_io_config),
    .io_in_0(Muxn_10_io_in_0),
    .io_in_1(Muxn_10_io_in_1),
    .io_in_2(Muxn_10_io_in_2),
    .io_in_3(Muxn_10_io_in_3),
    .io_in_4(Muxn_10_io_in_4),
    .io_out(Muxn_10_io_out)
  );
  Muxn_147 Muxn_11 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_11_io_config),
    .io_in_0(Muxn_11_io_in_0),
    .io_in_1(Muxn_11_io_in_1),
    .io_in_2(Muxn_11_io_in_2),
    .io_in_3(Muxn_11_io_in_3),
    .io_in_4(Muxn_11_io_in_4),
    .io_out(Muxn_11_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNE_0 = Muxn_2_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinNE_1 = Muxn_3_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinSE_0 = Muxn_4_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSE_1 = Muxn_5_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSW_0 = Muxn_6_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_ipinSW_1 = Muxn_7_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_otrackW_0 = _T_12; // @[Interconnect.scala 430:21 Interconnect.scala 477:45]
  assign io_otrackN_0 = _T_14; // @[Interconnect.scala 431:21 Interconnect.scala 477:45]
  assign io_otrackE_0 = _T_16; // @[Interconnect.scala 432:21 Interconnect.scala 477:45]
  assign io_otrackS_0 = _T_18; // @[Interconnect.scala 433:21 Interconnect.scala 477:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 464:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 466:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 483:23]
  assign Muxn_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 483:23]
  assign Muxn_1_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 483:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 483:23]
  assign Muxn_3_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 483:23]
  assign Muxn_4_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 483:23]
  assign Muxn_5_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[13:12]; // @[Interconnect.scala 483:23]
  assign Muxn_6_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[15:14]; // @[Interconnect.scala 483:23]
  assign Muxn_7_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[18:16]; // @[Interconnect.scala 483:23]
  assign Muxn_8_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[21:19]; // @[Interconnect.scala 483:23]
  assign Muxn_9_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_config = ConfigMem_io_out_0[24:22]; // @[Interconnect.scala 483:23]
  assign Muxn_10_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_config = ConfigMem_io_out_0[27:25]; // @[Interconnect.scala 483:23]
  assign Muxn_11_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_4 = io_itrackE_0; // @[Interconnect.scala 475:63]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_12 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  _T_14 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  _T_16 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  _T_18 = _RAND_3[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_12 <= Muxn_8_io_out;
    _T_14 <= Muxn_9_io_out;
    _T_16 <= Muxn_10_io_out;
    _T_18 <= Muxn_11_io_out;
  end
endmodule
module GIB_52(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
  wire  ConfigMem_clock; // @[Interconnect.scala 463:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 463:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 463:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 463:21]
  wire [27:0] ConfigMem_io_out_0; // @[Interconnect.scala 463:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_6_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_7_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_10_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_11_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_out; // @[Interconnect.scala 473:25]
  wire  _T_1 = 10'h74 == io_cfg_addr[11:2]; // @[Interconnect.scala 464:50]
  ConfigMem_90 ConfigMem ( // @[Interconnect.scala 463:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_148 Muxn ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_out(Muxn_io_out)
  );
  Muxn_148 Muxn_1 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_out(Muxn_1_io_out)
  );
  Muxn_148 Muxn_2 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_in_3(Muxn_2_io_in_3),
    .io_out(Muxn_2_io_out)
  );
  Muxn_148 Muxn_3 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_in_3(Muxn_3_io_in_3),
    .io_out(Muxn_3_io_out)
  );
  Muxn_148 Muxn_4 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_in_3(Muxn_4_io_in_3),
    .io_out(Muxn_4_io_out)
  );
  Muxn_148 Muxn_5 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_in_3(Muxn_5_io_in_3),
    .io_out(Muxn_5_io_out)
  );
  Muxn_148 Muxn_6 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_out(Muxn_6_io_out)
  );
  Muxn_148 Muxn_7 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_out(Muxn_7_io_out)
  );
  Muxn_147 Muxn_8 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_147 Muxn_9 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  Muxn_147 Muxn_10 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_10_io_config),
    .io_in_0(Muxn_10_io_in_0),
    .io_in_1(Muxn_10_io_in_1),
    .io_in_2(Muxn_10_io_in_2),
    .io_in_3(Muxn_10_io_in_3),
    .io_in_4(Muxn_10_io_in_4),
    .io_out(Muxn_10_io_out)
  );
  Muxn_147 Muxn_11 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_11_io_config),
    .io_in_0(Muxn_11_io_in_0),
    .io_in_1(Muxn_11_io_in_1),
    .io_in_2(Muxn_11_io_in_2),
    .io_in_3(Muxn_11_io_in_3),
    .io_in_4(Muxn_11_io_in_4),
    .io_out(Muxn_11_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNE_0 = Muxn_2_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinNE_1 = Muxn_3_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinSE_0 = Muxn_4_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSE_1 = Muxn_5_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSW_0 = Muxn_6_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_ipinSW_1 = Muxn_7_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_otrackW_0 = Muxn_8_io_out; // @[Interconnect.scala 430:21 Interconnect.scala 479:45]
  assign io_otrackN_0 = Muxn_9_io_out; // @[Interconnect.scala 431:21 Interconnect.scala 479:45]
  assign io_otrackE_0 = Muxn_10_io_out; // @[Interconnect.scala 432:21 Interconnect.scala 479:45]
  assign io_otrackS_0 = Muxn_11_io_out; // @[Interconnect.scala 433:21 Interconnect.scala 479:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 464:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 466:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 483:23]
  assign Muxn_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 483:23]
  assign Muxn_1_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 483:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 483:23]
  assign Muxn_3_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 483:23]
  assign Muxn_4_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 483:23]
  assign Muxn_5_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[13:12]; // @[Interconnect.scala 483:23]
  assign Muxn_6_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[15:14]; // @[Interconnect.scala 483:23]
  assign Muxn_7_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[18:16]; // @[Interconnect.scala 483:23]
  assign Muxn_8_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[21:19]; // @[Interconnect.scala 483:23]
  assign Muxn_9_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_config = ConfigMem_io_out_0[24:22]; // @[Interconnect.scala 483:23]
  assign Muxn_10_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_config = ConfigMem_io_out_0[27:25]; // @[Interconnect.scala 483:23]
  assign Muxn_11_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_4 = io_itrackE_0; // @[Interconnect.scala 475:63]
endmodule
module GIB_53(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire  ConfigMem_clock; // @[Interconnect.scala 463:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 463:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 463:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 463:21]
  wire [14:0] ConfigMem_io_out_0; // @[Interconnect.scala 463:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 473:25]
  wire  Muxn_2_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 473:25]
  wire  Muxn_3_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_6_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_7_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 473:25]
  wire  _T_1 = 10'h75 == io_cfg_addr[11:2]; // @[Interconnect.scala 464:50]
  reg [31:0] _T_8; // @[Interconnect.scala 477:55]
  reg [31:0] _T_10; // @[Interconnect.scala 477:55]
  reg [31:0] _T_14; // @[Interconnect.scala 477:55]
  ConfigMem_89 ConfigMem ( // @[Interconnect.scala 463:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_145 Muxn ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_out(Muxn_io_out)
  );
  Muxn_145 Muxn_1 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_out(Muxn_1_io_out)
  );
  Muxn Muxn_2 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_out(Muxn_2_io_out)
  );
  Muxn Muxn_3 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_out(Muxn_3_io_out)
  );
  Muxn_145 Muxn_4 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_out(Muxn_4_io_out)
  );
  Muxn_148 Muxn_5 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_in_3(Muxn_5_io_in_3),
    .io_out(Muxn_5_io_out)
  );
  Muxn_147 Muxn_6 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_in_4(Muxn_6_io_in_4),
    .io_out(Muxn_6_io_out)
  );
  Muxn_148 Muxn_7 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_out(Muxn_7_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinSW_0 = Muxn_2_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_ipinSW_1 = Muxn_3_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_otrackW_0 = _T_8; // @[Interconnect.scala 430:21 Interconnect.scala 477:45]
  assign io_otrackN_0 = _T_10; // @[Interconnect.scala 431:21 Interconnect.scala 477:45]
  assign io_otrackS_0 = _T_14; // @[Interconnect.scala 433:21 Interconnect.scala 477:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 464:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 466:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 483:23]
  assign Muxn_io_in_0 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_1 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_2 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 483:23]
  assign Muxn_1_io_in_0 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_1 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_2 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[4]; // @[Interconnect.scala 483:23]
  assign Muxn_2_io_in_0 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_1 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[5]; // @[Interconnect.scala 483:23]
  assign Muxn_3_io_in_0 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_1 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 483:23]
  assign Muxn_4_io_in_0 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_1 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_2 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 483:23]
  assign Muxn_5_io_in_0 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_1 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_2 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[12:10]; // @[Interconnect.scala 483:23]
  assign Muxn_6_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[14:13]; // @[Interconnect.scala 483:23]
  assign Muxn_7_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_1 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_3 = 32'h0; // @[Interconnect.scala 475:63]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_8 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  _T_10 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  _T_14 = _RAND_2[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_8 <= Muxn_4_io_out;
    _T_10 <= Muxn_5_io_out;
    _T_14 <= Muxn_7_io_out;
  end
endmodule
module GIB_54(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
  wire  ConfigMem_clock; // @[Interconnect.scala 463:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 463:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 463:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 463:21]
  wire [14:0] ConfigMem_io_out_0; // @[Interconnect.scala 463:21]
  wire  Muxn_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 473:25]
  wire  Muxn_1_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_4_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_6_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_7_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 473:25]
  wire  _T_1 = 10'h7f == io_cfg_addr[11:2]; // @[Interconnect.scala 464:50]
  ConfigMem_89 ConfigMem ( // @[Interconnect.scala 463:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn Muxn ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_out(Muxn_io_out)
  );
  Muxn Muxn_1 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_out(Muxn_1_io_out)
  );
  Muxn_145 Muxn_2 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_out(Muxn_2_io_out)
  );
  Muxn_145 Muxn_3 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_out(Muxn_3_io_out)
  );
  Muxn_147 Muxn_4 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_in_3(Muxn_4_io_in_3),
    .io_in_4(Muxn_4_io_in_4),
    .io_out(Muxn_4_io_out)
  );
  Muxn_148 Muxn_5 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_in_3(Muxn_5_io_in_3),
    .io_out(Muxn_5_io_out)
  );
  Muxn_145 Muxn_6 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_out(Muxn_6_io_out)
  );
  Muxn_148 Muxn_7 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_out(Muxn_7_io_out)
  );
  assign io_ipinNE_0 = Muxn_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinNE_1 = Muxn_1_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinSE_0 = Muxn_2_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSE_1 = Muxn_3_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_otrackN_0 = Muxn_5_io_out; // @[Interconnect.scala 431:21 Interconnect.scala 479:45]
  assign io_otrackE_0 = Muxn_6_io_out; // @[Interconnect.scala 432:21 Interconnect.scala 479:45]
  assign io_otrackS_0 = Muxn_7_io_out; // @[Interconnect.scala 433:21 Interconnect.scala 479:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 464:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 466:21]
  assign Muxn_io_config = ConfigMem_io_out_0[0]; // @[Interconnect.scala 483:23]
  assign Muxn_io_in_0 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_1 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[1]; // @[Interconnect.scala 483:23]
  assign Muxn_1_io_in_0 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_1 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 483:23]
  assign Muxn_2_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_1 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 483:23]
  assign Muxn_3_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_1 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[8:6]; // @[Interconnect.scala 483:23]
  assign Muxn_4_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[10:9]; // @[Interconnect.scala 483:23]
  assign Muxn_5_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_1 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[12:11]; // @[Interconnect.scala 483:23]
  assign Muxn_6_io_in_0 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_1 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_2 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[14:13]; // @[Interconnect.scala 483:23]
  assign Muxn_7_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_1 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
endmodule
module GIB_55(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire  ConfigMem_clock; // @[Interconnect.scala 463:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 463:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 463:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 463:21]
  wire [27:0] ConfigMem_io_out_0; // @[Interconnect.scala 463:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_6_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_7_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_10_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_11_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_out; // @[Interconnect.scala 473:25]
  wire  _T_1 = 10'h80 == io_cfg_addr[11:2]; // @[Interconnect.scala 464:50]
  reg [31:0] _T_12; // @[Interconnect.scala 477:55]
  reg [31:0] _T_14; // @[Interconnect.scala 477:55]
  reg [31:0] _T_16; // @[Interconnect.scala 477:55]
  reg [31:0] _T_18; // @[Interconnect.scala 477:55]
  ConfigMem_90 ConfigMem ( // @[Interconnect.scala 463:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_148 Muxn ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_out(Muxn_io_out)
  );
  Muxn_148 Muxn_1 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_out(Muxn_1_io_out)
  );
  Muxn_148 Muxn_2 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_in_3(Muxn_2_io_in_3),
    .io_out(Muxn_2_io_out)
  );
  Muxn_148 Muxn_3 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_in_3(Muxn_3_io_in_3),
    .io_out(Muxn_3_io_out)
  );
  Muxn_148 Muxn_4 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_in_3(Muxn_4_io_in_3),
    .io_out(Muxn_4_io_out)
  );
  Muxn_148 Muxn_5 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_in_3(Muxn_5_io_in_3),
    .io_out(Muxn_5_io_out)
  );
  Muxn_148 Muxn_6 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_out(Muxn_6_io_out)
  );
  Muxn_148 Muxn_7 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_out(Muxn_7_io_out)
  );
  Muxn_147 Muxn_8 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_147 Muxn_9 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  Muxn_147 Muxn_10 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_10_io_config),
    .io_in_0(Muxn_10_io_in_0),
    .io_in_1(Muxn_10_io_in_1),
    .io_in_2(Muxn_10_io_in_2),
    .io_in_3(Muxn_10_io_in_3),
    .io_in_4(Muxn_10_io_in_4),
    .io_out(Muxn_10_io_out)
  );
  Muxn_147 Muxn_11 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_11_io_config),
    .io_in_0(Muxn_11_io_in_0),
    .io_in_1(Muxn_11_io_in_1),
    .io_in_2(Muxn_11_io_in_2),
    .io_in_3(Muxn_11_io_in_3),
    .io_in_4(Muxn_11_io_in_4),
    .io_out(Muxn_11_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNE_0 = Muxn_2_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinNE_1 = Muxn_3_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinSE_0 = Muxn_4_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSE_1 = Muxn_5_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSW_0 = Muxn_6_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_ipinSW_1 = Muxn_7_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_otrackW_0 = _T_12; // @[Interconnect.scala 430:21 Interconnect.scala 477:45]
  assign io_otrackN_0 = _T_14; // @[Interconnect.scala 431:21 Interconnect.scala 477:45]
  assign io_otrackE_0 = _T_16; // @[Interconnect.scala 432:21 Interconnect.scala 477:45]
  assign io_otrackS_0 = _T_18; // @[Interconnect.scala 433:21 Interconnect.scala 477:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 464:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 466:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 483:23]
  assign Muxn_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 483:23]
  assign Muxn_1_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 483:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 483:23]
  assign Muxn_3_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 483:23]
  assign Muxn_4_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 483:23]
  assign Muxn_5_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[13:12]; // @[Interconnect.scala 483:23]
  assign Muxn_6_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[15:14]; // @[Interconnect.scala 483:23]
  assign Muxn_7_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[18:16]; // @[Interconnect.scala 483:23]
  assign Muxn_8_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[21:19]; // @[Interconnect.scala 483:23]
  assign Muxn_9_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_config = ConfigMem_io_out_0[24:22]; // @[Interconnect.scala 483:23]
  assign Muxn_10_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_config = ConfigMem_io_out_0[27:25]; // @[Interconnect.scala 483:23]
  assign Muxn_11_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_4 = io_itrackE_0; // @[Interconnect.scala 475:63]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_12 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  _T_14 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  _T_16 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  _T_18 = _RAND_3[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_12 <= Muxn_8_io_out;
    _T_14 <= Muxn_9_io_out;
    _T_16 <= Muxn_10_io_out;
    _T_18 <= Muxn_11_io_out;
  end
endmodule
module GIB_56(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
  wire  ConfigMem_clock; // @[Interconnect.scala 463:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 463:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 463:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 463:21]
  wire [27:0] ConfigMem_io_out_0; // @[Interconnect.scala 463:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_6_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_7_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_10_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_11_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_out; // @[Interconnect.scala 473:25]
  wire  _T_1 = 10'h81 == io_cfg_addr[11:2]; // @[Interconnect.scala 464:50]
  ConfigMem_90 ConfigMem ( // @[Interconnect.scala 463:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_148 Muxn ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_out(Muxn_io_out)
  );
  Muxn_148 Muxn_1 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_out(Muxn_1_io_out)
  );
  Muxn_148 Muxn_2 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_in_3(Muxn_2_io_in_3),
    .io_out(Muxn_2_io_out)
  );
  Muxn_148 Muxn_3 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_in_3(Muxn_3_io_in_3),
    .io_out(Muxn_3_io_out)
  );
  Muxn_148 Muxn_4 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_in_3(Muxn_4_io_in_3),
    .io_out(Muxn_4_io_out)
  );
  Muxn_148 Muxn_5 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_in_3(Muxn_5_io_in_3),
    .io_out(Muxn_5_io_out)
  );
  Muxn_148 Muxn_6 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_out(Muxn_6_io_out)
  );
  Muxn_148 Muxn_7 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_out(Muxn_7_io_out)
  );
  Muxn_147 Muxn_8 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_147 Muxn_9 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  Muxn_147 Muxn_10 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_10_io_config),
    .io_in_0(Muxn_10_io_in_0),
    .io_in_1(Muxn_10_io_in_1),
    .io_in_2(Muxn_10_io_in_2),
    .io_in_3(Muxn_10_io_in_3),
    .io_in_4(Muxn_10_io_in_4),
    .io_out(Muxn_10_io_out)
  );
  Muxn_147 Muxn_11 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_11_io_config),
    .io_in_0(Muxn_11_io_in_0),
    .io_in_1(Muxn_11_io_in_1),
    .io_in_2(Muxn_11_io_in_2),
    .io_in_3(Muxn_11_io_in_3),
    .io_in_4(Muxn_11_io_in_4),
    .io_out(Muxn_11_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNE_0 = Muxn_2_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinNE_1 = Muxn_3_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinSE_0 = Muxn_4_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSE_1 = Muxn_5_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSW_0 = Muxn_6_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_ipinSW_1 = Muxn_7_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_otrackW_0 = Muxn_8_io_out; // @[Interconnect.scala 430:21 Interconnect.scala 479:45]
  assign io_otrackN_0 = Muxn_9_io_out; // @[Interconnect.scala 431:21 Interconnect.scala 479:45]
  assign io_otrackE_0 = Muxn_10_io_out; // @[Interconnect.scala 432:21 Interconnect.scala 479:45]
  assign io_otrackS_0 = Muxn_11_io_out; // @[Interconnect.scala 433:21 Interconnect.scala 479:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 464:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 466:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 483:23]
  assign Muxn_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 483:23]
  assign Muxn_1_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 483:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 483:23]
  assign Muxn_3_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 483:23]
  assign Muxn_4_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 483:23]
  assign Muxn_5_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[13:12]; // @[Interconnect.scala 483:23]
  assign Muxn_6_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[15:14]; // @[Interconnect.scala 483:23]
  assign Muxn_7_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[18:16]; // @[Interconnect.scala 483:23]
  assign Muxn_8_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[21:19]; // @[Interconnect.scala 483:23]
  assign Muxn_9_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_config = ConfigMem_io_out_0[24:22]; // @[Interconnect.scala 483:23]
  assign Muxn_10_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_config = ConfigMem_io_out_0[27:25]; // @[Interconnect.scala 483:23]
  assign Muxn_11_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_4 = io_itrackE_0; // @[Interconnect.scala 475:63]
endmodule
module GIB_57(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire  ConfigMem_clock; // @[Interconnect.scala 463:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 463:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 463:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 463:21]
  wire [27:0] ConfigMem_io_out_0; // @[Interconnect.scala 463:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_6_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_7_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_10_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_11_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_out; // @[Interconnect.scala 473:25]
  wire  _T_1 = 10'h82 == io_cfg_addr[11:2]; // @[Interconnect.scala 464:50]
  reg [31:0] _T_12; // @[Interconnect.scala 477:55]
  reg [31:0] _T_14; // @[Interconnect.scala 477:55]
  reg [31:0] _T_16; // @[Interconnect.scala 477:55]
  reg [31:0] _T_18; // @[Interconnect.scala 477:55]
  ConfigMem_90 ConfigMem ( // @[Interconnect.scala 463:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_148 Muxn ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_out(Muxn_io_out)
  );
  Muxn_148 Muxn_1 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_out(Muxn_1_io_out)
  );
  Muxn_148 Muxn_2 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_in_3(Muxn_2_io_in_3),
    .io_out(Muxn_2_io_out)
  );
  Muxn_148 Muxn_3 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_in_3(Muxn_3_io_in_3),
    .io_out(Muxn_3_io_out)
  );
  Muxn_148 Muxn_4 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_in_3(Muxn_4_io_in_3),
    .io_out(Muxn_4_io_out)
  );
  Muxn_148 Muxn_5 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_in_3(Muxn_5_io_in_3),
    .io_out(Muxn_5_io_out)
  );
  Muxn_148 Muxn_6 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_out(Muxn_6_io_out)
  );
  Muxn_148 Muxn_7 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_out(Muxn_7_io_out)
  );
  Muxn_147 Muxn_8 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_147 Muxn_9 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  Muxn_147 Muxn_10 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_10_io_config),
    .io_in_0(Muxn_10_io_in_0),
    .io_in_1(Muxn_10_io_in_1),
    .io_in_2(Muxn_10_io_in_2),
    .io_in_3(Muxn_10_io_in_3),
    .io_in_4(Muxn_10_io_in_4),
    .io_out(Muxn_10_io_out)
  );
  Muxn_147 Muxn_11 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_11_io_config),
    .io_in_0(Muxn_11_io_in_0),
    .io_in_1(Muxn_11_io_in_1),
    .io_in_2(Muxn_11_io_in_2),
    .io_in_3(Muxn_11_io_in_3),
    .io_in_4(Muxn_11_io_in_4),
    .io_out(Muxn_11_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNE_0 = Muxn_2_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinNE_1 = Muxn_3_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinSE_0 = Muxn_4_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSE_1 = Muxn_5_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSW_0 = Muxn_6_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_ipinSW_1 = Muxn_7_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_otrackW_0 = _T_12; // @[Interconnect.scala 430:21 Interconnect.scala 477:45]
  assign io_otrackN_0 = _T_14; // @[Interconnect.scala 431:21 Interconnect.scala 477:45]
  assign io_otrackE_0 = _T_16; // @[Interconnect.scala 432:21 Interconnect.scala 477:45]
  assign io_otrackS_0 = _T_18; // @[Interconnect.scala 433:21 Interconnect.scala 477:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 464:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 466:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 483:23]
  assign Muxn_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 483:23]
  assign Muxn_1_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 483:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 483:23]
  assign Muxn_3_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 483:23]
  assign Muxn_4_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 483:23]
  assign Muxn_5_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[13:12]; // @[Interconnect.scala 483:23]
  assign Muxn_6_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[15:14]; // @[Interconnect.scala 483:23]
  assign Muxn_7_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[18:16]; // @[Interconnect.scala 483:23]
  assign Muxn_8_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[21:19]; // @[Interconnect.scala 483:23]
  assign Muxn_9_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_config = ConfigMem_io_out_0[24:22]; // @[Interconnect.scala 483:23]
  assign Muxn_10_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_config = ConfigMem_io_out_0[27:25]; // @[Interconnect.scala 483:23]
  assign Muxn_11_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_4 = io_itrackE_0; // @[Interconnect.scala 475:63]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_12 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  _T_14 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  _T_16 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  _T_18 = _RAND_3[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_12 <= Muxn_8_io_out;
    _T_14 <= Muxn_9_io_out;
    _T_16 <= Muxn_10_io_out;
    _T_18 <= Muxn_11_io_out;
  end
endmodule
module GIB_58(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
  wire  ConfigMem_clock; // @[Interconnect.scala 463:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 463:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 463:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 463:21]
  wire [27:0] ConfigMem_io_out_0; // @[Interconnect.scala 463:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_6_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_7_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_10_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_11_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_out; // @[Interconnect.scala 473:25]
  wire  _T_1 = 10'h83 == io_cfg_addr[11:2]; // @[Interconnect.scala 464:50]
  ConfigMem_90 ConfigMem ( // @[Interconnect.scala 463:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_148 Muxn ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_out(Muxn_io_out)
  );
  Muxn_148 Muxn_1 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_out(Muxn_1_io_out)
  );
  Muxn_148 Muxn_2 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_in_3(Muxn_2_io_in_3),
    .io_out(Muxn_2_io_out)
  );
  Muxn_148 Muxn_3 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_in_3(Muxn_3_io_in_3),
    .io_out(Muxn_3_io_out)
  );
  Muxn_148 Muxn_4 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_in_3(Muxn_4_io_in_3),
    .io_out(Muxn_4_io_out)
  );
  Muxn_148 Muxn_5 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_in_3(Muxn_5_io_in_3),
    .io_out(Muxn_5_io_out)
  );
  Muxn_148 Muxn_6 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_out(Muxn_6_io_out)
  );
  Muxn_148 Muxn_7 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_out(Muxn_7_io_out)
  );
  Muxn_147 Muxn_8 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_147 Muxn_9 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  Muxn_147 Muxn_10 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_10_io_config),
    .io_in_0(Muxn_10_io_in_0),
    .io_in_1(Muxn_10_io_in_1),
    .io_in_2(Muxn_10_io_in_2),
    .io_in_3(Muxn_10_io_in_3),
    .io_in_4(Muxn_10_io_in_4),
    .io_out(Muxn_10_io_out)
  );
  Muxn_147 Muxn_11 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_11_io_config),
    .io_in_0(Muxn_11_io_in_0),
    .io_in_1(Muxn_11_io_in_1),
    .io_in_2(Muxn_11_io_in_2),
    .io_in_3(Muxn_11_io_in_3),
    .io_in_4(Muxn_11_io_in_4),
    .io_out(Muxn_11_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNE_0 = Muxn_2_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinNE_1 = Muxn_3_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinSE_0 = Muxn_4_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSE_1 = Muxn_5_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSW_0 = Muxn_6_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_ipinSW_1 = Muxn_7_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_otrackW_0 = Muxn_8_io_out; // @[Interconnect.scala 430:21 Interconnect.scala 479:45]
  assign io_otrackN_0 = Muxn_9_io_out; // @[Interconnect.scala 431:21 Interconnect.scala 479:45]
  assign io_otrackE_0 = Muxn_10_io_out; // @[Interconnect.scala 432:21 Interconnect.scala 479:45]
  assign io_otrackS_0 = Muxn_11_io_out; // @[Interconnect.scala 433:21 Interconnect.scala 479:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 464:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 466:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 483:23]
  assign Muxn_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 483:23]
  assign Muxn_1_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 483:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 483:23]
  assign Muxn_3_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 483:23]
  assign Muxn_4_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 483:23]
  assign Muxn_5_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[13:12]; // @[Interconnect.scala 483:23]
  assign Muxn_6_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[15:14]; // @[Interconnect.scala 483:23]
  assign Muxn_7_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[18:16]; // @[Interconnect.scala 483:23]
  assign Muxn_8_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[21:19]; // @[Interconnect.scala 483:23]
  assign Muxn_9_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_config = ConfigMem_io_out_0[24:22]; // @[Interconnect.scala 483:23]
  assign Muxn_10_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_config = ConfigMem_io_out_0[27:25]; // @[Interconnect.scala 483:23]
  assign Muxn_11_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_4 = io_itrackE_0; // @[Interconnect.scala 475:63]
endmodule
module GIB_59(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire  ConfigMem_clock; // @[Interconnect.scala 463:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 463:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 463:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 463:21]
  wire [27:0] ConfigMem_io_out_0; // @[Interconnect.scala 463:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_6_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_7_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_10_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_11_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_out; // @[Interconnect.scala 473:25]
  wire  _T_1 = 10'h84 == io_cfg_addr[11:2]; // @[Interconnect.scala 464:50]
  reg [31:0] _T_12; // @[Interconnect.scala 477:55]
  reg [31:0] _T_14; // @[Interconnect.scala 477:55]
  reg [31:0] _T_16; // @[Interconnect.scala 477:55]
  reg [31:0] _T_18; // @[Interconnect.scala 477:55]
  ConfigMem_90 ConfigMem ( // @[Interconnect.scala 463:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_148 Muxn ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_out(Muxn_io_out)
  );
  Muxn_148 Muxn_1 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_out(Muxn_1_io_out)
  );
  Muxn_148 Muxn_2 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_in_3(Muxn_2_io_in_3),
    .io_out(Muxn_2_io_out)
  );
  Muxn_148 Muxn_3 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_in_3(Muxn_3_io_in_3),
    .io_out(Muxn_3_io_out)
  );
  Muxn_148 Muxn_4 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_in_3(Muxn_4_io_in_3),
    .io_out(Muxn_4_io_out)
  );
  Muxn_148 Muxn_5 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_in_3(Muxn_5_io_in_3),
    .io_out(Muxn_5_io_out)
  );
  Muxn_148 Muxn_6 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_out(Muxn_6_io_out)
  );
  Muxn_148 Muxn_7 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_out(Muxn_7_io_out)
  );
  Muxn_147 Muxn_8 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_147 Muxn_9 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  Muxn_147 Muxn_10 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_10_io_config),
    .io_in_0(Muxn_10_io_in_0),
    .io_in_1(Muxn_10_io_in_1),
    .io_in_2(Muxn_10_io_in_2),
    .io_in_3(Muxn_10_io_in_3),
    .io_in_4(Muxn_10_io_in_4),
    .io_out(Muxn_10_io_out)
  );
  Muxn_147 Muxn_11 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_11_io_config),
    .io_in_0(Muxn_11_io_in_0),
    .io_in_1(Muxn_11_io_in_1),
    .io_in_2(Muxn_11_io_in_2),
    .io_in_3(Muxn_11_io_in_3),
    .io_in_4(Muxn_11_io_in_4),
    .io_out(Muxn_11_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNE_0 = Muxn_2_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinNE_1 = Muxn_3_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinSE_0 = Muxn_4_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSE_1 = Muxn_5_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSW_0 = Muxn_6_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_ipinSW_1 = Muxn_7_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_otrackW_0 = _T_12; // @[Interconnect.scala 430:21 Interconnect.scala 477:45]
  assign io_otrackN_0 = _T_14; // @[Interconnect.scala 431:21 Interconnect.scala 477:45]
  assign io_otrackE_0 = _T_16; // @[Interconnect.scala 432:21 Interconnect.scala 477:45]
  assign io_otrackS_0 = _T_18; // @[Interconnect.scala 433:21 Interconnect.scala 477:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 464:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 466:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 483:23]
  assign Muxn_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 483:23]
  assign Muxn_1_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 483:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 483:23]
  assign Muxn_3_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 483:23]
  assign Muxn_4_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 483:23]
  assign Muxn_5_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[13:12]; // @[Interconnect.scala 483:23]
  assign Muxn_6_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[15:14]; // @[Interconnect.scala 483:23]
  assign Muxn_7_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[18:16]; // @[Interconnect.scala 483:23]
  assign Muxn_8_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[21:19]; // @[Interconnect.scala 483:23]
  assign Muxn_9_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_config = ConfigMem_io_out_0[24:22]; // @[Interconnect.scala 483:23]
  assign Muxn_10_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_config = ConfigMem_io_out_0[27:25]; // @[Interconnect.scala 483:23]
  assign Muxn_11_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_4 = io_itrackE_0; // @[Interconnect.scala 475:63]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_12 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  _T_14 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  _T_16 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  _T_18 = _RAND_3[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_12 <= Muxn_8_io_out;
    _T_14 <= Muxn_9_io_out;
    _T_16 <= Muxn_10_io_out;
    _T_18 <= Muxn_11_io_out;
  end
endmodule
module GIB_60(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
  wire  ConfigMem_clock; // @[Interconnect.scala 463:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 463:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 463:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 463:21]
  wire [27:0] ConfigMem_io_out_0; // @[Interconnect.scala 463:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_6_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_7_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_10_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_11_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_out; // @[Interconnect.scala 473:25]
  wire  _T_1 = 10'h85 == io_cfg_addr[11:2]; // @[Interconnect.scala 464:50]
  ConfigMem_90 ConfigMem ( // @[Interconnect.scala 463:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_148 Muxn ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_out(Muxn_io_out)
  );
  Muxn_148 Muxn_1 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_out(Muxn_1_io_out)
  );
  Muxn_148 Muxn_2 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_in_3(Muxn_2_io_in_3),
    .io_out(Muxn_2_io_out)
  );
  Muxn_148 Muxn_3 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_in_3(Muxn_3_io_in_3),
    .io_out(Muxn_3_io_out)
  );
  Muxn_148 Muxn_4 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_in_3(Muxn_4_io_in_3),
    .io_out(Muxn_4_io_out)
  );
  Muxn_148 Muxn_5 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_in_3(Muxn_5_io_in_3),
    .io_out(Muxn_5_io_out)
  );
  Muxn_148 Muxn_6 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_out(Muxn_6_io_out)
  );
  Muxn_148 Muxn_7 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_out(Muxn_7_io_out)
  );
  Muxn_147 Muxn_8 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_147 Muxn_9 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  Muxn_147 Muxn_10 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_10_io_config),
    .io_in_0(Muxn_10_io_in_0),
    .io_in_1(Muxn_10_io_in_1),
    .io_in_2(Muxn_10_io_in_2),
    .io_in_3(Muxn_10_io_in_3),
    .io_in_4(Muxn_10_io_in_4),
    .io_out(Muxn_10_io_out)
  );
  Muxn_147 Muxn_11 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_11_io_config),
    .io_in_0(Muxn_11_io_in_0),
    .io_in_1(Muxn_11_io_in_1),
    .io_in_2(Muxn_11_io_in_2),
    .io_in_3(Muxn_11_io_in_3),
    .io_in_4(Muxn_11_io_in_4),
    .io_out(Muxn_11_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNE_0 = Muxn_2_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinNE_1 = Muxn_3_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinSE_0 = Muxn_4_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSE_1 = Muxn_5_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSW_0 = Muxn_6_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_ipinSW_1 = Muxn_7_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_otrackW_0 = Muxn_8_io_out; // @[Interconnect.scala 430:21 Interconnect.scala 479:45]
  assign io_otrackN_0 = Muxn_9_io_out; // @[Interconnect.scala 431:21 Interconnect.scala 479:45]
  assign io_otrackE_0 = Muxn_10_io_out; // @[Interconnect.scala 432:21 Interconnect.scala 479:45]
  assign io_otrackS_0 = Muxn_11_io_out; // @[Interconnect.scala 433:21 Interconnect.scala 479:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 464:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 466:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 483:23]
  assign Muxn_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 483:23]
  assign Muxn_1_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 483:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 483:23]
  assign Muxn_3_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 483:23]
  assign Muxn_4_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 483:23]
  assign Muxn_5_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[13:12]; // @[Interconnect.scala 483:23]
  assign Muxn_6_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[15:14]; // @[Interconnect.scala 483:23]
  assign Muxn_7_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[18:16]; // @[Interconnect.scala 483:23]
  assign Muxn_8_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[21:19]; // @[Interconnect.scala 483:23]
  assign Muxn_9_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_config = ConfigMem_io_out_0[24:22]; // @[Interconnect.scala 483:23]
  assign Muxn_10_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_config = ConfigMem_io_out_0[27:25]; // @[Interconnect.scala 483:23]
  assign Muxn_11_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_4 = io_itrackE_0; // @[Interconnect.scala 475:63]
endmodule
module GIB_61(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire  ConfigMem_clock; // @[Interconnect.scala 463:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 463:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 463:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 463:21]
  wire [27:0] ConfigMem_io_out_0; // @[Interconnect.scala 463:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_6_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_7_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_10_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_11_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_out; // @[Interconnect.scala 473:25]
  wire  _T_1 = 10'h86 == io_cfg_addr[11:2]; // @[Interconnect.scala 464:50]
  reg [31:0] _T_12; // @[Interconnect.scala 477:55]
  reg [31:0] _T_14; // @[Interconnect.scala 477:55]
  reg [31:0] _T_16; // @[Interconnect.scala 477:55]
  reg [31:0] _T_18; // @[Interconnect.scala 477:55]
  ConfigMem_90 ConfigMem ( // @[Interconnect.scala 463:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_148 Muxn ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_out(Muxn_io_out)
  );
  Muxn_148 Muxn_1 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_out(Muxn_1_io_out)
  );
  Muxn_148 Muxn_2 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_in_3(Muxn_2_io_in_3),
    .io_out(Muxn_2_io_out)
  );
  Muxn_148 Muxn_3 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_in_3(Muxn_3_io_in_3),
    .io_out(Muxn_3_io_out)
  );
  Muxn_148 Muxn_4 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_in_3(Muxn_4_io_in_3),
    .io_out(Muxn_4_io_out)
  );
  Muxn_148 Muxn_5 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_in_3(Muxn_5_io_in_3),
    .io_out(Muxn_5_io_out)
  );
  Muxn_148 Muxn_6 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_out(Muxn_6_io_out)
  );
  Muxn_148 Muxn_7 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_out(Muxn_7_io_out)
  );
  Muxn_147 Muxn_8 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_147 Muxn_9 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  Muxn_147 Muxn_10 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_10_io_config),
    .io_in_0(Muxn_10_io_in_0),
    .io_in_1(Muxn_10_io_in_1),
    .io_in_2(Muxn_10_io_in_2),
    .io_in_3(Muxn_10_io_in_3),
    .io_in_4(Muxn_10_io_in_4),
    .io_out(Muxn_10_io_out)
  );
  Muxn_147 Muxn_11 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_11_io_config),
    .io_in_0(Muxn_11_io_in_0),
    .io_in_1(Muxn_11_io_in_1),
    .io_in_2(Muxn_11_io_in_2),
    .io_in_3(Muxn_11_io_in_3),
    .io_in_4(Muxn_11_io_in_4),
    .io_out(Muxn_11_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNE_0 = Muxn_2_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinNE_1 = Muxn_3_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinSE_0 = Muxn_4_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSE_1 = Muxn_5_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSW_0 = Muxn_6_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_ipinSW_1 = Muxn_7_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_otrackW_0 = _T_12; // @[Interconnect.scala 430:21 Interconnect.scala 477:45]
  assign io_otrackN_0 = _T_14; // @[Interconnect.scala 431:21 Interconnect.scala 477:45]
  assign io_otrackE_0 = _T_16; // @[Interconnect.scala 432:21 Interconnect.scala 477:45]
  assign io_otrackS_0 = _T_18; // @[Interconnect.scala 433:21 Interconnect.scala 477:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 464:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 466:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 483:23]
  assign Muxn_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 483:23]
  assign Muxn_1_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 483:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 483:23]
  assign Muxn_3_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 483:23]
  assign Muxn_4_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 483:23]
  assign Muxn_5_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[13:12]; // @[Interconnect.scala 483:23]
  assign Muxn_6_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[15:14]; // @[Interconnect.scala 483:23]
  assign Muxn_7_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[18:16]; // @[Interconnect.scala 483:23]
  assign Muxn_8_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[21:19]; // @[Interconnect.scala 483:23]
  assign Muxn_9_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_config = ConfigMem_io_out_0[24:22]; // @[Interconnect.scala 483:23]
  assign Muxn_10_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_config = ConfigMem_io_out_0[27:25]; // @[Interconnect.scala 483:23]
  assign Muxn_11_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_4 = io_itrackE_0; // @[Interconnect.scala 475:63]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_12 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  _T_14 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  _T_16 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  _T_18 = _RAND_3[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_12 <= Muxn_8_io_out;
    _T_14 <= Muxn_9_io_out;
    _T_16 <= Muxn_10_io_out;
    _T_18 <= Muxn_11_io_out;
  end
endmodule
module GIB_62(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
  wire  ConfigMem_clock; // @[Interconnect.scala 463:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 463:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 463:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 463:21]
  wire [14:0] ConfigMem_io_out_0; // @[Interconnect.scala 463:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 473:25]
  wire  Muxn_2_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 473:25]
  wire  Muxn_3_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_6_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_7_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 473:25]
  wire  _T_1 = 10'h87 == io_cfg_addr[11:2]; // @[Interconnect.scala 464:50]
  ConfigMem_89 ConfigMem ( // @[Interconnect.scala 463:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_145 Muxn ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_out(Muxn_io_out)
  );
  Muxn_145 Muxn_1 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_out(Muxn_1_io_out)
  );
  Muxn Muxn_2 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_out(Muxn_2_io_out)
  );
  Muxn Muxn_3 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_out(Muxn_3_io_out)
  );
  Muxn_145 Muxn_4 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_out(Muxn_4_io_out)
  );
  Muxn_148 Muxn_5 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_in_3(Muxn_5_io_in_3),
    .io_out(Muxn_5_io_out)
  );
  Muxn_147 Muxn_6 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_in_4(Muxn_6_io_in_4),
    .io_out(Muxn_6_io_out)
  );
  Muxn_148 Muxn_7 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_out(Muxn_7_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinSW_0 = Muxn_2_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_ipinSW_1 = Muxn_3_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_otrackW_0 = Muxn_4_io_out; // @[Interconnect.scala 430:21 Interconnect.scala 479:45]
  assign io_otrackN_0 = Muxn_5_io_out; // @[Interconnect.scala 431:21 Interconnect.scala 479:45]
  assign io_otrackS_0 = Muxn_7_io_out; // @[Interconnect.scala 433:21 Interconnect.scala 479:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 464:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 466:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 483:23]
  assign Muxn_io_in_0 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_1 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_2 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 483:23]
  assign Muxn_1_io_in_0 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_1 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_2 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[4]; // @[Interconnect.scala 483:23]
  assign Muxn_2_io_in_0 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_1 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[5]; // @[Interconnect.scala 483:23]
  assign Muxn_3_io_in_0 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_1 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 483:23]
  assign Muxn_4_io_in_0 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_1 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_2 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 483:23]
  assign Muxn_5_io_in_0 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_1 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_2 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[12:10]; // @[Interconnect.scala 483:23]
  assign Muxn_6_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[14:13]; // @[Interconnect.scala 483:23]
  assign Muxn_7_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_1 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_3 = 32'h0; // @[Interconnect.scala 475:63]
endmodule
module GIB_63(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire  ConfigMem_clock; // @[Interconnect.scala 463:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 463:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 463:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 463:21]
  wire [14:0] ConfigMem_io_out_0; // @[Interconnect.scala 463:21]
  wire  Muxn_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 473:25]
  wire  Muxn_1_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_4_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_6_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_7_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 473:25]
  wire  _T_1 = 10'h91 == io_cfg_addr[11:2]; // @[Interconnect.scala 464:50]
  reg [31:0] _T_10; // @[Interconnect.scala 477:55]
  reg [31:0] _T_12; // @[Interconnect.scala 477:55]
  reg [31:0] _T_14; // @[Interconnect.scala 477:55]
  ConfigMem_89 ConfigMem ( // @[Interconnect.scala 463:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn Muxn ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_out(Muxn_io_out)
  );
  Muxn Muxn_1 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_out(Muxn_1_io_out)
  );
  Muxn_145 Muxn_2 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_out(Muxn_2_io_out)
  );
  Muxn_145 Muxn_3 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_out(Muxn_3_io_out)
  );
  Muxn_147 Muxn_4 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_in_3(Muxn_4_io_in_3),
    .io_in_4(Muxn_4_io_in_4),
    .io_out(Muxn_4_io_out)
  );
  Muxn_148 Muxn_5 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_in_3(Muxn_5_io_in_3),
    .io_out(Muxn_5_io_out)
  );
  Muxn_145 Muxn_6 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_out(Muxn_6_io_out)
  );
  Muxn_148 Muxn_7 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_out(Muxn_7_io_out)
  );
  assign io_ipinNE_0 = Muxn_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinNE_1 = Muxn_1_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinSE_0 = Muxn_2_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSE_1 = Muxn_3_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_otrackN_0 = _T_10; // @[Interconnect.scala 431:21 Interconnect.scala 477:45]
  assign io_otrackE_0 = _T_12; // @[Interconnect.scala 432:21 Interconnect.scala 477:45]
  assign io_otrackS_0 = _T_14; // @[Interconnect.scala 433:21 Interconnect.scala 477:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 464:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 466:21]
  assign Muxn_io_config = ConfigMem_io_out_0[0]; // @[Interconnect.scala 483:23]
  assign Muxn_io_in_0 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_1 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[1]; // @[Interconnect.scala 483:23]
  assign Muxn_1_io_in_0 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_1 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 483:23]
  assign Muxn_2_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_1 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 483:23]
  assign Muxn_3_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_1 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[8:6]; // @[Interconnect.scala 483:23]
  assign Muxn_4_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[10:9]; // @[Interconnect.scala 483:23]
  assign Muxn_5_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_1 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[12:11]; // @[Interconnect.scala 483:23]
  assign Muxn_6_io_in_0 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_1 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_2 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[14:13]; // @[Interconnect.scala 483:23]
  assign Muxn_7_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_1 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_10 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  _T_12 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  _T_14 = _RAND_2[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_10 <= Muxn_5_io_out;
    _T_12 <= Muxn_6_io_out;
    _T_14 <= Muxn_7_io_out;
  end
endmodule
module GIB_64(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
  wire  ConfigMem_clock; // @[Interconnect.scala 463:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 463:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 463:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 463:21]
  wire [27:0] ConfigMem_io_out_0; // @[Interconnect.scala 463:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_6_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_7_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_10_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_11_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_out; // @[Interconnect.scala 473:25]
  wire  _T_1 = 10'h92 == io_cfg_addr[11:2]; // @[Interconnect.scala 464:50]
  ConfigMem_90 ConfigMem ( // @[Interconnect.scala 463:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_148 Muxn ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_out(Muxn_io_out)
  );
  Muxn_148 Muxn_1 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_out(Muxn_1_io_out)
  );
  Muxn_148 Muxn_2 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_in_3(Muxn_2_io_in_3),
    .io_out(Muxn_2_io_out)
  );
  Muxn_148 Muxn_3 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_in_3(Muxn_3_io_in_3),
    .io_out(Muxn_3_io_out)
  );
  Muxn_148 Muxn_4 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_in_3(Muxn_4_io_in_3),
    .io_out(Muxn_4_io_out)
  );
  Muxn_148 Muxn_5 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_in_3(Muxn_5_io_in_3),
    .io_out(Muxn_5_io_out)
  );
  Muxn_148 Muxn_6 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_out(Muxn_6_io_out)
  );
  Muxn_148 Muxn_7 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_out(Muxn_7_io_out)
  );
  Muxn_147 Muxn_8 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_147 Muxn_9 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  Muxn_147 Muxn_10 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_10_io_config),
    .io_in_0(Muxn_10_io_in_0),
    .io_in_1(Muxn_10_io_in_1),
    .io_in_2(Muxn_10_io_in_2),
    .io_in_3(Muxn_10_io_in_3),
    .io_in_4(Muxn_10_io_in_4),
    .io_out(Muxn_10_io_out)
  );
  Muxn_147 Muxn_11 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_11_io_config),
    .io_in_0(Muxn_11_io_in_0),
    .io_in_1(Muxn_11_io_in_1),
    .io_in_2(Muxn_11_io_in_2),
    .io_in_3(Muxn_11_io_in_3),
    .io_in_4(Muxn_11_io_in_4),
    .io_out(Muxn_11_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNE_0 = Muxn_2_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinNE_1 = Muxn_3_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinSE_0 = Muxn_4_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSE_1 = Muxn_5_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSW_0 = Muxn_6_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_ipinSW_1 = Muxn_7_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_otrackW_0 = Muxn_8_io_out; // @[Interconnect.scala 430:21 Interconnect.scala 479:45]
  assign io_otrackN_0 = Muxn_9_io_out; // @[Interconnect.scala 431:21 Interconnect.scala 479:45]
  assign io_otrackE_0 = Muxn_10_io_out; // @[Interconnect.scala 432:21 Interconnect.scala 479:45]
  assign io_otrackS_0 = Muxn_11_io_out; // @[Interconnect.scala 433:21 Interconnect.scala 479:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 464:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 466:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 483:23]
  assign Muxn_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 483:23]
  assign Muxn_1_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 483:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 483:23]
  assign Muxn_3_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 483:23]
  assign Muxn_4_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 483:23]
  assign Muxn_5_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[13:12]; // @[Interconnect.scala 483:23]
  assign Muxn_6_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[15:14]; // @[Interconnect.scala 483:23]
  assign Muxn_7_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[18:16]; // @[Interconnect.scala 483:23]
  assign Muxn_8_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[21:19]; // @[Interconnect.scala 483:23]
  assign Muxn_9_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_config = ConfigMem_io_out_0[24:22]; // @[Interconnect.scala 483:23]
  assign Muxn_10_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_config = ConfigMem_io_out_0[27:25]; // @[Interconnect.scala 483:23]
  assign Muxn_11_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_4 = io_itrackE_0; // @[Interconnect.scala 475:63]
endmodule
module GIB_65(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire  ConfigMem_clock; // @[Interconnect.scala 463:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 463:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 463:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 463:21]
  wire [27:0] ConfigMem_io_out_0; // @[Interconnect.scala 463:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_6_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_7_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_10_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_11_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_out; // @[Interconnect.scala 473:25]
  wire  _T_1 = 10'h93 == io_cfg_addr[11:2]; // @[Interconnect.scala 464:50]
  reg [31:0] _T_12; // @[Interconnect.scala 477:55]
  reg [31:0] _T_14; // @[Interconnect.scala 477:55]
  reg [31:0] _T_16; // @[Interconnect.scala 477:55]
  reg [31:0] _T_18; // @[Interconnect.scala 477:55]
  ConfigMem_90 ConfigMem ( // @[Interconnect.scala 463:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_148 Muxn ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_out(Muxn_io_out)
  );
  Muxn_148 Muxn_1 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_out(Muxn_1_io_out)
  );
  Muxn_148 Muxn_2 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_in_3(Muxn_2_io_in_3),
    .io_out(Muxn_2_io_out)
  );
  Muxn_148 Muxn_3 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_in_3(Muxn_3_io_in_3),
    .io_out(Muxn_3_io_out)
  );
  Muxn_148 Muxn_4 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_in_3(Muxn_4_io_in_3),
    .io_out(Muxn_4_io_out)
  );
  Muxn_148 Muxn_5 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_in_3(Muxn_5_io_in_3),
    .io_out(Muxn_5_io_out)
  );
  Muxn_148 Muxn_6 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_out(Muxn_6_io_out)
  );
  Muxn_148 Muxn_7 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_out(Muxn_7_io_out)
  );
  Muxn_147 Muxn_8 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_147 Muxn_9 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  Muxn_147 Muxn_10 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_10_io_config),
    .io_in_0(Muxn_10_io_in_0),
    .io_in_1(Muxn_10_io_in_1),
    .io_in_2(Muxn_10_io_in_2),
    .io_in_3(Muxn_10_io_in_3),
    .io_in_4(Muxn_10_io_in_4),
    .io_out(Muxn_10_io_out)
  );
  Muxn_147 Muxn_11 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_11_io_config),
    .io_in_0(Muxn_11_io_in_0),
    .io_in_1(Muxn_11_io_in_1),
    .io_in_2(Muxn_11_io_in_2),
    .io_in_3(Muxn_11_io_in_3),
    .io_in_4(Muxn_11_io_in_4),
    .io_out(Muxn_11_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNE_0 = Muxn_2_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinNE_1 = Muxn_3_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinSE_0 = Muxn_4_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSE_1 = Muxn_5_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSW_0 = Muxn_6_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_ipinSW_1 = Muxn_7_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_otrackW_0 = _T_12; // @[Interconnect.scala 430:21 Interconnect.scala 477:45]
  assign io_otrackN_0 = _T_14; // @[Interconnect.scala 431:21 Interconnect.scala 477:45]
  assign io_otrackE_0 = _T_16; // @[Interconnect.scala 432:21 Interconnect.scala 477:45]
  assign io_otrackS_0 = _T_18; // @[Interconnect.scala 433:21 Interconnect.scala 477:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 464:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 466:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 483:23]
  assign Muxn_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 483:23]
  assign Muxn_1_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 483:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 483:23]
  assign Muxn_3_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 483:23]
  assign Muxn_4_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 483:23]
  assign Muxn_5_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[13:12]; // @[Interconnect.scala 483:23]
  assign Muxn_6_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[15:14]; // @[Interconnect.scala 483:23]
  assign Muxn_7_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[18:16]; // @[Interconnect.scala 483:23]
  assign Muxn_8_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[21:19]; // @[Interconnect.scala 483:23]
  assign Muxn_9_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_config = ConfigMem_io_out_0[24:22]; // @[Interconnect.scala 483:23]
  assign Muxn_10_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_config = ConfigMem_io_out_0[27:25]; // @[Interconnect.scala 483:23]
  assign Muxn_11_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_4 = io_itrackE_0; // @[Interconnect.scala 475:63]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_12 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  _T_14 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  _T_16 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  _T_18 = _RAND_3[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_12 <= Muxn_8_io_out;
    _T_14 <= Muxn_9_io_out;
    _T_16 <= Muxn_10_io_out;
    _T_18 <= Muxn_11_io_out;
  end
endmodule
module GIB_66(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
  wire  ConfigMem_clock; // @[Interconnect.scala 463:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 463:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 463:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 463:21]
  wire [27:0] ConfigMem_io_out_0; // @[Interconnect.scala 463:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_6_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_7_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_10_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_11_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_out; // @[Interconnect.scala 473:25]
  wire  _T_1 = 10'h94 == io_cfg_addr[11:2]; // @[Interconnect.scala 464:50]
  ConfigMem_90 ConfigMem ( // @[Interconnect.scala 463:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_148 Muxn ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_out(Muxn_io_out)
  );
  Muxn_148 Muxn_1 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_out(Muxn_1_io_out)
  );
  Muxn_148 Muxn_2 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_in_3(Muxn_2_io_in_3),
    .io_out(Muxn_2_io_out)
  );
  Muxn_148 Muxn_3 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_in_3(Muxn_3_io_in_3),
    .io_out(Muxn_3_io_out)
  );
  Muxn_148 Muxn_4 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_in_3(Muxn_4_io_in_3),
    .io_out(Muxn_4_io_out)
  );
  Muxn_148 Muxn_5 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_in_3(Muxn_5_io_in_3),
    .io_out(Muxn_5_io_out)
  );
  Muxn_148 Muxn_6 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_out(Muxn_6_io_out)
  );
  Muxn_148 Muxn_7 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_out(Muxn_7_io_out)
  );
  Muxn_147 Muxn_8 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_147 Muxn_9 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  Muxn_147 Muxn_10 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_10_io_config),
    .io_in_0(Muxn_10_io_in_0),
    .io_in_1(Muxn_10_io_in_1),
    .io_in_2(Muxn_10_io_in_2),
    .io_in_3(Muxn_10_io_in_3),
    .io_in_4(Muxn_10_io_in_4),
    .io_out(Muxn_10_io_out)
  );
  Muxn_147 Muxn_11 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_11_io_config),
    .io_in_0(Muxn_11_io_in_0),
    .io_in_1(Muxn_11_io_in_1),
    .io_in_2(Muxn_11_io_in_2),
    .io_in_3(Muxn_11_io_in_3),
    .io_in_4(Muxn_11_io_in_4),
    .io_out(Muxn_11_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNE_0 = Muxn_2_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinNE_1 = Muxn_3_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinSE_0 = Muxn_4_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSE_1 = Muxn_5_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSW_0 = Muxn_6_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_ipinSW_1 = Muxn_7_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_otrackW_0 = Muxn_8_io_out; // @[Interconnect.scala 430:21 Interconnect.scala 479:45]
  assign io_otrackN_0 = Muxn_9_io_out; // @[Interconnect.scala 431:21 Interconnect.scala 479:45]
  assign io_otrackE_0 = Muxn_10_io_out; // @[Interconnect.scala 432:21 Interconnect.scala 479:45]
  assign io_otrackS_0 = Muxn_11_io_out; // @[Interconnect.scala 433:21 Interconnect.scala 479:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 464:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 466:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 483:23]
  assign Muxn_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 483:23]
  assign Muxn_1_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 483:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 483:23]
  assign Muxn_3_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 483:23]
  assign Muxn_4_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 483:23]
  assign Muxn_5_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[13:12]; // @[Interconnect.scala 483:23]
  assign Muxn_6_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[15:14]; // @[Interconnect.scala 483:23]
  assign Muxn_7_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[18:16]; // @[Interconnect.scala 483:23]
  assign Muxn_8_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[21:19]; // @[Interconnect.scala 483:23]
  assign Muxn_9_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_config = ConfigMem_io_out_0[24:22]; // @[Interconnect.scala 483:23]
  assign Muxn_10_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_config = ConfigMem_io_out_0[27:25]; // @[Interconnect.scala 483:23]
  assign Muxn_11_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_4 = io_itrackE_0; // @[Interconnect.scala 475:63]
endmodule
module GIB_67(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire  ConfigMem_clock; // @[Interconnect.scala 463:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 463:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 463:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 463:21]
  wire [27:0] ConfigMem_io_out_0; // @[Interconnect.scala 463:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_6_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_7_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_10_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_11_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_out; // @[Interconnect.scala 473:25]
  wire  _T_1 = 10'h95 == io_cfg_addr[11:2]; // @[Interconnect.scala 464:50]
  reg [31:0] _T_12; // @[Interconnect.scala 477:55]
  reg [31:0] _T_14; // @[Interconnect.scala 477:55]
  reg [31:0] _T_16; // @[Interconnect.scala 477:55]
  reg [31:0] _T_18; // @[Interconnect.scala 477:55]
  ConfigMem_90 ConfigMem ( // @[Interconnect.scala 463:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_148 Muxn ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_out(Muxn_io_out)
  );
  Muxn_148 Muxn_1 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_out(Muxn_1_io_out)
  );
  Muxn_148 Muxn_2 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_in_3(Muxn_2_io_in_3),
    .io_out(Muxn_2_io_out)
  );
  Muxn_148 Muxn_3 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_in_3(Muxn_3_io_in_3),
    .io_out(Muxn_3_io_out)
  );
  Muxn_148 Muxn_4 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_in_3(Muxn_4_io_in_3),
    .io_out(Muxn_4_io_out)
  );
  Muxn_148 Muxn_5 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_in_3(Muxn_5_io_in_3),
    .io_out(Muxn_5_io_out)
  );
  Muxn_148 Muxn_6 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_out(Muxn_6_io_out)
  );
  Muxn_148 Muxn_7 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_out(Muxn_7_io_out)
  );
  Muxn_147 Muxn_8 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_147 Muxn_9 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  Muxn_147 Muxn_10 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_10_io_config),
    .io_in_0(Muxn_10_io_in_0),
    .io_in_1(Muxn_10_io_in_1),
    .io_in_2(Muxn_10_io_in_2),
    .io_in_3(Muxn_10_io_in_3),
    .io_in_4(Muxn_10_io_in_4),
    .io_out(Muxn_10_io_out)
  );
  Muxn_147 Muxn_11 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_11_io_config),
    .io_in_0(Muxn_11_io_in_0),
    .io_in_1(Muxn_11_io_in_1),
    .io_in_2(Muxn_11_io_in_2),
    .io_in_3(Muxn_11_io_in_3),
    .io_in_4(Muxn_11_io_in_4),
    .io_out(Muxn_11_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNE_0 = Muxn_2_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinNE_1 = Muxn_3_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinSE_0 = Muxn_4_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSE_1 = Muxn_5_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSW_0 = Muxn_6_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_ipinSW_1 = Muxn_7_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_otrackW_0 = _T_12; // @[Interconnect.scala 430:21 Interconnect.scala 477:45]
  assign io_otrackN_0 = _T_14; // @[Interconnect.scala 431:21 Interconnect.scala 477:45]
  assign io_otrackE_0 = _T_16; // @[Interconnect.scala 432:21 Interconnect.scala 477:45]
  assign io_otrackS_0 = _T_18; // @[Interconnect.scala 433:21 Interconnect.scala 477:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 464:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 466:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 483:23]
  assign Muxn_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 483:23]
  assign Muxn_1_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 483:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 483:23]
  assign Muxn_3_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 483:23]
  assign Muxn_4_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 483:23]
  assign Muxn_5_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[13:12]; // @[Interconnect.scala 483:23]
  assign Muxn_6_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[15:14]; // @[Interconnect.scala 483:23]
  assign Muxn_7_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[18:16]; // @[Interconnect.scala 483:23]
  assign Muxn_8_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[21:19]; // @[Interconnect.scala 483:23]
  assign Muxn_9_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_config = ConfigMem_io_out_0[24:22]; // @[Interconnect.scala 483:23]
  assign Muxn_10_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_config = ConfigMem_io_out_0[27:25]; // @[Interconnect.scala 483:23]
  assign Muxn_11_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_4 = io_itrackE_0; // @[Interconnect.scala 475:63]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_12 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  _T_14 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  _T_16 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  _T_18 = _RAND_3[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_12 <= Muxn_8_io_out;
    _T_14 <= Muxn_9_io_out;
    _T_16 <= Muxn_10_io_out;
    _T_18 <= Muxn_11_io_out;
  end
endmodule
module GIB_68(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
  wire  ConfigMem_clock; // @[Interconnect.scala 463:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 463:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 463:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 463:21]
  wire [27:0] ConfigMem_io_out_0; // @[Interconnect.scala 463:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_6_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_7_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_10_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_11_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_out; // @[Interconnect.scala 473:25]
  wire  _T_1 = 10'h96 == io_cfg_addr[11:2]; // @[Interconnect.scala 464:50]
  ConfigMem_90 ConfigMem ( // @[Interconnect.scala 463:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_148 Muxn ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_out(Muxn_io_out)
  );
  Muxn_148 Muxn_1 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_out(Muxn_1_io_out)
  );
  Muxn_148 Muxn_2 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_in_3(Muxn_2_io_in_3),
    .io_out(Muxn_2_io_out)
  );
  Muxn_148 Muxn_3 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_in_3(Muxn_3_io_in_3),
    .io_out(Muxn_3_io_out)
  );
  Muxn_148 Muxn_4 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_in_3(Muxn_4_io_in_3),
    .io_out(Muxn_4_io_out)
  );
  Muxn_148 Muxn_5 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_in_3(Muxn_5_io_in_3),
    .io_out(Muxn_5_io_out)
  );
  Muxn_148 Muxn_6 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_out(Muxn_6_io_out)
  );
  Muxn_148 Muxn_7 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_out(Muxn_7_io_out)
  );
  Muxn_147 Muxn_8 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_147 Muxn_9 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  Muxn_147 Muxn_10 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_10_io_config),
    .io_in_0(Muxn_10_io_in_0),
    .io_in_1(Muxn_10_io_in_1),
    .io_in_2(Muxn_10_io_in_2),
    .io_in_3(Muxn_10_io_in_3),
    .io_in_4(Muxn_10_io_in_4),
    .io_out(Muxn_10_io_out)
  );
  Muxn_147 Muxn_11 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_11_io_config),
    .io_in_0(Muxn_11_io_in_0),
    .io_in_1(Muxn_11_io_in_1),
    .io_in_2(Muxn_11_io_in_2),
    .io_in_3(Muxn_11_io_in_3),
    .io_in_4(Muxn_11_io_in_4),
    .io_out(Muxn_11_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNE_0 = Muxn_2_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinNE_1 = Muxn_3_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinSE_0 = Muxn_4_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSE_1 = Muxn_5_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSW_0 = Muxn_6_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_ipinSW_1 = Muxn_7_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_otrackW_0 = Muxn_8_io_out; // @[Interconnect.scala 430:21 Interconnect.scala 479:45]
  assign io_otrackN_0 = Muxn_9_io_out; // @[Interconnect.scala 431:21 Interconnect.scala 479:45]
  assign io_otrackE_0 = Muxn_10_io_out; // @[Interconnect.scala 432:21 Interconnect.scala 479:45]
  assign io_otrackS_0 = Muxn_11_io_out; // @[Interconnect.scala 433:21 Interconnect.scala 479:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 464:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 466:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 483:23]
  assign Muxn_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 483:23]
  assign Muxn_1_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 483:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 483:23]
  assign Muxn_3_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 483:23]
  assign Muxn_4_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 483:23]
  assign Muxn_5_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[13:12]; // @[Interconnect.scala 483:23]
  assign Muxn_6_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[15:14]; // @[Interconnect.scala 483:23]
  assign Muxn_7_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[18:16]; // @[Interconnect.scala 483:23]
  assign Muxn_8_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[21:19]; // @[Interconnect.scala 483:23]
  assign Muxn_9_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_config = ConfigMem_io_out_0[24:22]; // @[Interconnect.scala 483:23]
  assign Muxn_10_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_config = ConfigMem_io_out_0[27:25]; // @[Interconnect.scala 483:23]
  assign Muxn_11_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_4 = io_itrackE_0; // @[Interconnect.scala 475:63]
endmodule
module GIB_69(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire  ConfigMem_clock; // @[Interconnect.scala 463:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 463:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 463:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 463:21]
  wire [27:0] ConfigMem_io_out_0; // @[Interconnect.scala 463:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_6_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_7_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_10_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_11_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_out; // @[Interconnect.scala 473:25]
  wire  _T_1 = 10'h97 == io_cfg_addr[11:2]; // @[Interconnect.scala 464:50]
  reg [31:0] _T_12; // @[Interconnect.scala 477:55]
  reg [31:0] _T_14; // @[Interconnect.scala 477:55]
  reg [31:0] _T_16; // @[Interconnect.scala 477:55]
  reg [31:0] _T_18; // @[Interconnect.scala 477:55]
  ConfigMem_90 ConfigMem ( // @[Interconnect.scala 463:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_148 Muxn ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_out(Muxn_io_out)
  );
  Muxn_148 Muxn_1 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_out(Muxn_1_io_out)
  );
  Muxn_148 Muxn_2 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_in_3(Muxn_2_io_in_3),
    .io_out(Muxn_2_io_out)
  );
  Muxn_148 Muxn_3 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_in_3(Muxn_3_io_in_3),
    .io_out(Muxn_3_io_out)
  );
  Muxn_148 Muxn_4 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_in_3(Muxn_4_io_in_3),
    .io_out(Muxn_4_io_out)
  );
  Muxn_148 Muxn_5 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_in_3(Muxn_5_io_in_3),
    .io_out(Muxn_5_io_out)
  );
  Muxn_148 Muxn_6 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_out(Muxn_6_io_out)
  );
  Muxn_148 Muxn_7 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_out(Muxn_7_io_out)
  );
  Muxn_147 Muxn_8 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_147 Muxn_9 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  Muxn_147 Muxn_10 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_10_io_config),
    .io_in_0(Muxn_10_io_in_0),
    .io_in_1(Muxn_10_io_in_1),
    .io_in_2(Muxn_10_io_in_2),
    .io_in_3(Muxn_10_io_in_3),
    .io_in_4(Muxn_10_io_in_4),
    .io_out(Muxn_10_io_out)
  );
  Muxn_147 Muxn_11 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_11_io_config),
    .io_in_0(Muxn_11_io_in_0),
    .io_in_1(Muxn_11_io_in_1),
    .io_in_2(Muxn_11_io_in_2),
    .io_in_3(Muxn_11_io_in_3),
    .io_in_4(Muxn_11_io_in_4),
    .io_out(Muxn_11_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNE_0 = Muxn_2_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinNE_1 = Muxn_3_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinSE_0 = Muxn_4_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSE_1 = Muxn_5_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSW_0 = Muxn_6_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_ipinSW_1 = Muxn_7_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_otrackW_0 = _T_12; // @[Interconnect.scala 430:21 Interconnect.scala 477:45]
  assign io_otrackN_0 = _T_14; // @[Interconnect.scala 431:21 Interconnect.scala 477:45]
  assign io_otrackE_0 = _T_16; // @[Interconnect.scala 432:21 Interconnect.scala 477:45]
  assign io_otrackS_0 = _T_18; // @[Interconnect.scala 433:21 Interconnect.scala 477:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 464:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 466:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 483:23]
  assign Muxn_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 483:23]
  assign Muxn_1_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 483:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 483:23]
  assign Muxn_3_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 483:23]
  assign Muxn_4_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 483:23]
  assign Muxn_5_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[13:12]; // @[Interconnect.scala 483:23]
  assign Muxn_6_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[15:14]; // @[Interconnect.scala 483:23]
  assign Muxn_7_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[18:16]; // @[Interconnect.scala 483:23]
  assign Muxn_8_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[21:19]; // @[Interconnect.scala 483:23]
  assign Muxn_9_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_config = ConfigMem_io_out_0[24:22]; // @[Interconnect.scala 483:23]
  assign Muxn_10_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_config = ConfigMem_io_out_0[27:25]; // @[Interconnect.scala 483:23]
  assign Muxn_11_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_4 = io_itrackE_0; // @[Interconnect.scala 475:63]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_12 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  _T_14 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  _T_16 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  _T_18 = _RAND_3[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_12 <= Muxn_8_io_out;
    _T_14 <= Muxn_9_io_out;
    _T_16 <= Muxn_10_io_out;
    _T_18 <= Muxn_11_io_out;
  end
endmodule
module GIB_70(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
  wire  ConfigMem_clock; // @[Interconnect.scala 463:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 463:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 463:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 463:21]
  wire [27:0] ConfigMem_io_out_0; // @[Interconnect.scala 463:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_6_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_7_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_10_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_10_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_11_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_11_io_out; // @[Interconnect.scala 473:25]
  wire  _T_1 = 10'h98 == io_cfg_addr[11:2]; // @[Interconnect.scala 464:50]
  ConfigMem_90 ConfigMem ( // @[Interconnect.scala 463:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_148 Muxn ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_out(Muxn_io_out)
  );
  Muxn_148 Muxn_1 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_out(Muxn_1_io_out)
  );
  Muxn_148 Muxn_2 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_in_3(Muxn_2_io_in_3),
    .io_out(Muxn_2_io_out)
  );
  Muxn_148 Muxn_3 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_in_3(Muxn_3_io_in_3),
    .io_out(Muxn_3_io_out)
  );
  Muxn_148 Muxn_4 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_in_3(Muxn_4_io_in_3),
    .io_out(Muxn_4_io_out)
  );
  Muxn_148 Muxn_5 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_in_3(Muxn_5_io_in_3),
    .io_out(Muxn_5_io_out)
  );
  Muxn_148 Muxn_6 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_out(Muxn_6_io_out)
  );
  Muxn_148 Muxn_7 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_out(Muxn_7_io_out)
  );
  Muxn_147 Muxn_8 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_147 Muxn_9 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  Muxn_147 Muxn_10 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_10_io_config),
    .io_in_0(Muxn_10_io_in_0),
    .io_in_1(Muxn_10_io_in_1),
    .io_in_2(Muxn_10_io_in_2),
    .io_in_3(Muxn_10_io_in_3),
    .io_in_4(Muxn_10_io_in_4),
    .io_out(Muxn_10_io_out)
  );
  Muxn_147 Muxn_11 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_11_io_config),
    .io_in_0(Muxn_11_io_in_0),
    .io_in_1(Muxn_11_io_in_1),
    .io_in_2(Muxn_11_io_in_2),
    .io_in_3(Muxn_11_io_in_3),
    .io_in_4(Muxn_11_io_in_4),
    .io_out(Muxn_11_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNE_0 = Muxn_2_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinNE_1 = Muxn_3_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinSE_0 = Muxn_4_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSE_1 = Muxn_5_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSW_0 = Muxn_6_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_ipinSW_1 = Muxn_7_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_otrackW_0 = Muxn_8_io_out; // @[Interconnect.scala 430:21 Interconnect.scala 479:45]
  assign io_otrackN_0 = Muxn_9_io_out; // @[Interconnect.scala 431:21 Interconnect.scala 479:45]
  assign io_otrackE_0 = Muxn_10_io_out; // @[Interconnect.scala 432:21 Interconnect.scala 479:45]
  assign io_otrackS_0 = Muxn_11_io_out; // @[Interconnect.scala 433:21 Interconnect.scala 479:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 464:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 466:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 483:23]
  assign Muxn_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 483:23]
  assign Muxn_1_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 483:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 483:23]
  assign Muxn_3_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 483:23]
  assign Muxn_4_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 483:23]
  assign Muxn_5_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[13:12]; // @[Interconnect.scala 483:23]
  assign Muxn_6_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[15:14]; // @[Interconnect.scala 483:23]
  assign Muxn_7_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[18:16]; // @[Interconnect.scala 483:23]
  assign Muxn_8_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[21:19]; // @[Interconnect.scala 483:23]
  assign Muxn_9_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_config = ConfigMem_io_out_0[24:22]; // @[Interconnect.scala 483:23]
  assign Muxn_10_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_10_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_config = ConfigMem_io_out_0[27:25]; // @[Interconnect.scala 483:23]
  assign Muxn_11_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_11_io_in_4 = io_itrackE_0; // @[Interconnect.scala 475:63]
endmodule
module GIB_71(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire  ConfigMem_clock; // @[Interconnect.scala 463:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 463:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 463:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 463:21]
  wire [14:0] ConfigMem_io_out_0; // @[Interconnect.scala 463:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 473:25]
  wire  Muxn_2_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 473:25]
  wire  Muxn_3_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_6_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_7_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 473:25]
  wire  _T_1 = 10'h99 == io_cfg_addr[11:2]; // @[Interconnect.scala 464:50]
  reg [31:0] _T_8; // @[Interconnect.scala 477:55]
  reg [31:0] _T_10; // @[Interconnect.scala 477:55]
  reg [31:0] _T_14; // @[Interconnect.scala 477:55]
  ConfigMem_89 ConfigMem ( // @[Interconnect.scala 463:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_145 Muxn ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_out(Muxn_io_out)
  );
  Muxn_145 Muxn_1 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_out(Muxn_1_io_out)
  );
  Muxn Muxn_2 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_out(Muxn_2_io_out)
  );
  Muxn Muxn_3 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_out(Muxn_3_io_out)
  );
  Muxn_145 Muxn_4 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_out(Muxn_4_io_out)
  );
  Muxn_148 Muxn_5 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_in_3(Muxn_5_io_in_3),
    .io_out(Muxn_5_io_out)
  );
  Muxn_147 Muxn_6 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_in_4(Muxn_6_io_in_4),
    .io_out(Muxn_6_io_out)
  );
  Muxn_148 Muxn_7 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_out(Muxn_7_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinSW_0 = Muxn_2_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_ipinSW_1 = Muxn_3_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_otrackW_0 = _T_8; // @[Interconnect.scala 430:21 Interconnect.scala 477:45]
  assign io_otrackN_0 = _T_10; // @[Interconnect.scala 431:21 Interconnect.scala 477:45]
  assign io_otrackS_0 = _T_14; // @[Interconnect.scala 433:21 Interconnect.scala 477:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 464:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 466:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 483:23]
  assign Muxn_io_in_0 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_1 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_2 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 483:23]
  assign Muxn_1_io_in_0 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_1 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_2 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[4]; // @[Interconnect.scala 483:23]
  assign Muxn_2_io_in_0 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_1 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[5]; // @[Interconnect.scala 483:23]
  assign Muxn_3_io_in_0 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_1 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 483:23]
  assign Muxn_4_io_in_0 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_1 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_2 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 483:23]
  assign Muxn_5_io_in_0 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_1 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_2 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_3 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[12:10]; // @[Interconnect.scala 483:23]
  assign Muxn_6_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_4 = io_itrackS_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[14:13]; // @[Interconnect.scala 483:23]
  assign Muxn_7_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_1 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_3 = 32'h0; // @[Interconnect.scala 475:63]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_8 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  _T_10 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  _T_14 = _RAND_2[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_8 <= Muxn_4_io_out;
    _T_10 <= Muxn_5_io_out;
    _T_14 <= Muxn_7_io_out;
  end
endmodule
module GIB_72(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  input  [31:0] io_opinSE_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0
);
  wire  ConfigMem_clock; // @[Interconnect.scala 463:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 463:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 463:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 463:21]
  wire [12:0] ConfigMem_io_out_0; // @[Interconnect.scala 463:21]
  wire  Muxn_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 473:25]
  wire  Muxn_1_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_3_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_6_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 473:25]
  wire  _T_1 = 10'ha3 == io_cfg_addr[11:2]; // @[Interconnect.scala 464:50]
  ConfigMem_88 ConfigMem ( // @[Interconnect.scala 463:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn Muxn ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_out(Muxn_io_out)
  );
  Muxn Muxn_1 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_out(Muxn_1_io_out)
  );
  Muxn_145 Muxn_2 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_out(Muxn_2_io_out)
  );
  Muxn_147 Muxn_3 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_in_3(Muxn_3_io_in_3),
    .io_in_4(Muxn_3_io_in_4),
    .io_out(Muxn_3_io_out)
  );
  Muxn_148 Muxn_4 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_in_3(Muxn_4_io_in_3),
    .io_out(Muxn_4_io_out)
  );
  Muxn_145 Muxn_5 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_out(Muxn_5_io_out)
  );
  Muxn_148 Muxn_6 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_out(Muxn_6_io_out)
  );
  assign io_ipinNE_0 = Muxn_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinNE_1 = Muxn_1_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinSE_0 = Muxn_2_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_otrackN_0 = Muxn_4_io_out; // @[Interconnect.scala 431:21 Interconnect.scala 479:45]
  assign io_otrackE_0 = Muxn_5_io_out; // @[Interconnect.scala 432:21 Interconnect.scala 479:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 464:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 466:21]
  assign Muxn_io_config = ConfigMem_io_out_0[0]; // @[Interconnect.scala 483:23]
  assign Muxn_io_in_0 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_1 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[1]; // @[Interconnect.scala 483:23]
  assign Muxn_1_io_in_0 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_1 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 483:23]
  assign Muxn_2_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_1 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[6:4]; // @[Interconnect.scala 483:23]
  assign Muxn_3_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_4 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[8:7]; // @[Interconnect.scala 483:23]
  assign Muxn_4_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_1 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_3 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[10:9]; // @[Interconnect.scala 483:23]
  assign Muxn_5_io_in_0 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_1 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_2 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[12:11]; // @[Interconnect.scala 483:23]
  assign Muxn_6_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_1 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
endmodule
module GIB_73(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire  ConfigMem_clock; // @[Interconnect.scala 463:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 463:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 463:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 463:21]
  wire [23:0] ConfigMem_io_out_0; // @[Interconnect.scala 463:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_6_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_7_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 473:25]
  wire  _T_1 = 10'ha4 == io_cfg_addr[11:2]; // @[Interconnect.scala 464:50]
  reg [31:0] _T_10; // @[Interconnect.scala 477:55]
  reg [31:0] _T_12; // @[Interconnect.scala 477:55]
  reg [31:0] _T_14; // @[Interconnect.scala 477:55]
  ConfigMem_81 ConfigMem ( // @[Interconnect.scala 463:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_148 Muxn ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_out(Muxn_io_out)
  );
  Muxn_148 Muxn_1 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_out(Muxn_1_io_out)
  );
  Muxn_148 Muxn_2 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_in_3(Muxn_2_io_in_3),
    .io_out(Muxn_2_io_out)
  );
  Muxn_148 Muxn_3 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_in_3(Muxn_3_io_in_3),
    .io_out(Muxn_3_io_out)
  );
  Muxn_148 Muxn_4 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_in_3(Muxn_4_io_in_3),
    .io_out(Muxn_4_io_out)
  );
  Muxn_148 Muxn_5 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_in_3(Muxn_5_io_in_3),
    .io_out(Muxn_5_io_out)
  );
  Muxn_147 Muxn_6 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_in_4(Muxn_6_io_in_4),
    .io_out(Muxn_6_io_out)
  );
  Muxn_147 Muxn_7 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_in_4(Muxn_7_io_in_4),
    .io_out(Muxn_7_io_out)
  );
  Muxn_147 Muxn_8 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_147 Muxn_9 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNE_0 = Muxn_2_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinNE_1 = Muxn_3_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinSE_0 = Muxn_4_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSW_0 = Muxn_5_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_otrackW_0 = _T_10; // @[Interconnect.scala 430:21 Interconnect.scala 477:45]
  assign io_otrackN_0 = _T_12; // @[Interconnect.scala 431:21 Interconnect.scala 477:45]
  assign io_otrackE_0 = _T_14; // @[Interconnect.scala 432:21 Interconnect.scala 477:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 464:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 466:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 483:23]
  assign Muxn_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_3 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 483:23]
  assign Muxn_1_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_3 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 483:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_3 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 483:23]
  assign Muxn_3_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_3 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 483:23]
  assign Muxn_4_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 483:23]
  assign Muxn_5_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[14:12]; // @[Interconnect.scala 483:23]
  assign Muxn_6_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_4 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[17:15]; // @[Interconnect.scala 483:23]
  assign Muxn_7_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_4 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[20:18]; // @[Interconnect.scala 483:23]
  assign Muxn_8_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_4 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[23:21]; // @[Interconnect.scala 483:23]
  assign Muxn_9_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_4 = io_itrackE_0; // @[Interconnect.scala 475:63]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_10 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  _T_12 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  _T_14 = _RAND_2[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_10 <= Muxn_6_io_out;
    _T_12 <= Muxn_7_io_out;
    _T_14 <= Muxn_8_io_out;
  end
endmodule
module GIB_74(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0
);
  wire  ConfigMem_clock; // @[Interconnect.scala 463:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 463:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 463:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 463:21]
  wire [23:0] ConfigMem_io_out_0; // @[Interconnect.scala 463:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_6_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_7_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 473:25]
  wire  _T_1 = 10'ha5 == io_cfg_addr[11:2]; // @[Interconnect.scala 464:50]
  ConfigMem_81 ConfigMem ( // @[Interconnect.scala 463:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_148 Muxn ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_out(Muxn_io_out)
  );
  Muxn_148 Muxn_1 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_out(Muxn_1_io_out)
  );
  Muxn_148 Muxn_2 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_in_3(Muxn_2_io_in_3),
    .io_out(Muxn_2_io_out)
  );
  Muxn_148 Muxn_3 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_in_3(Muxn_3_io_in_3),
    .io_out(Muxn_3_io_out)
  );
  Muxn_148 Muxn_4 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_in_3(Muxn_4_io_in_3),
    .io_out(Muxn_4_io_out)
  );
  Muxn_148 Muxn_5 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_in_3(Muxn_5_io_in_3),
    .io_out(Muxn_5_io_out)
  );
  Muxn_147 Muxn_6 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_in_4(Muxn_6_io_in_4),
    .io_out(Muxn_6_io_out)
  );
  Muxn_147 Muxn_7 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_in_4(Muxn_7_io_in_4),
    .io_out(Muxn_7_io_out)
  );
  Muxn_147 Muxn_8 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_147 Muxn_9 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNE_0 = Muxn_2_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinNE_1 = Muxn_3_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinSE_0 = Muxn_4_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSW_0 = Muxn_5_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_otrackW_0 = Muxn_6_io_out; // @[Interconnect.scala 430:21 Interconnect.scala 479:45]
  assign io_otrackN_0 = Muxn_7_io_out; // @[Interconnect.scala 431:21 Interconnect.scala 479:45]
  assign io_otrackE_0 = Muxn_8_io_out; // @[Interconnect.scala 432:21 Interconnect.scala 479:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 464:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 466:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 483:23]
  assign Muxn_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_3 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 483:23]
  assign Muxn_1_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_3 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 483:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_3 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 483:23]
  assign Muxn_3_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_3 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 483:23]
  assign Muxn_4_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 483:23]
  assign Muxn_5_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[14:12]; // @[Interconnect.scala 483:23]
  assign Muxn_6_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_4 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[17:15]; // @[Interconnect.scala 483:23]
  assign Muxn_7_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_4 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[20:18]; // @[Interconnect.scala 483:23]
  assign Muxn_8_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_4 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[23:21]; // @[Interconnect.scala 483:23]
  assign Muxn_9_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_4 = io_itrackE_0; // @[Interconnect.scala 475:63]
endmodule
module GIB_75(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire  ConfigMem_clock; // @[Interconnect.scala 463:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 463:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 463:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 463:21]
  wire [23:0] ConfigMem_io_out_0; // @[Interconnect.scala 463:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_6_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_7_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 473:25]
  wire  _T_1 = 10'ha6 == io_cfg_addr[11:2]; // @[Interconnect.scala 464:50]
  reg [31:0] _T_10; // @[Interconnect.scala 477:55]
  reg [31:0] _T_12; // @[Interconnect.scala 477:55]
  reg [31:0] _T_14; // @[Interconnect.scala 477:55]
  ConfigMem_81 ConfigMem ( // @[Interconnect.scala 463:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_148 Muxn ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_out(Muxn_io_out)
  );
  Muxn_148 Muxn_1 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_out(Muxn_1_io_out)
  );
  Muxn_148 Muxn_2 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_in_3(Muxn_2_io_in_3),
    .io_out(Muxn_2_io_out)
  );
  Muxn_148 Muxn_3 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_in_3(Muxn_3_io_in_3),
    .io_out(Muxn_3_io_out)
  );
  Muxn_148 Muxn_4 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_in_3(Muxn_4_io_in_3),
    .io_out(Muxn_4_io_out)
  );
  Muxn_148 Muxn_5 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_in_3(Muxn_5_io_in_3),
    .io_out(Muxn_5_io_out)
  );
  Muxn_147 Muxn_6 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_in_4(Muxn_6_io_in_4),
    .io_out(Muxn_6_io_out)
  );
  Muxn_147 Muxn_7 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_in_4(Muxn_7_io_in_4),
    .io_out(Muxn_7_io_out)
  );
  Muxn_147 Muxn_8 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_147 Muxn_9 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNE_0 = Muxn_2_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinNE_1 = Muxn_3_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinSE_0 = Muxn_4_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSW_0 = Muxn_5_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_otrackW_0 = _T_10; // @[Interconnect.scala 430:21 Interconnect.scala 477:45]
  assign io_otrackN_0 = _T_12; // @[Interconnect.scala 431:21 Interconnect.scala 477:45]
  assign io_otrackE_0 = _T_14; // @[Interconnect.scala 432:21 Interconnect.scala 477:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 464:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 466:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 483:23]
  assign Muxn_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_3 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 483:23]
  assign Muxn_1_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_3 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 483:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_3 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 483:23]
  assign Muxn_3_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_3 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 483:23]
  assign Muxn_4_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 483:23]
  assign Muxn_5_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[14:12]; // @[Interconnect.scala 483:23]
  assign Muxn_6_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_4 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[17:15]; // @[Interconnect.scala 483:23]
  assign Muxn_7_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_4 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[20:18]; // @[Interconnect.scala 483:23]
  assign Muxn_8_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_4 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[23:21]; // @[Interconnect.scala 483:23]
  assign Muxn_9_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_4 = io_itrackE_0; // @[Interconnect.scala 475:63]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_10 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  _T_12 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  _T_14 = _RAND_2[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_10 <= Muxn_6_io_out;
    _T_12 <= Muxn_7_io_out;
    _T_14 <= Muxn_8_io_out;
  end
endmodule
module GIB_76(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0
);
  wire  ConfigMem_clock; // @[Interconnect.scala 463:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 463:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 463:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 463:21]
  wire [23:0] ConfigMem_io_out_0; // @[Interconnect.scala 463:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_6_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_7_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 473:25]
  wire  _T_1 = 10'ha7 == io_cfg_addr[11:2]; // @[Interconnect.scala 464:50]
  ConfigMem_81 ConfigMem ( // @[Interconnect.scala 463:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_148 Muxn ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_out(Muxn_io_out)
  );
  Muxn_148 Muxn_1 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_out(Muxn_1_io_out)
  );
  Muxn_148 Muxn_2 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_in_3(Muxn_2_io_in_3),
    .io_out(Muxn_2_io_out)
  );
  Muxn_148 Muxn_3 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_in_3(Muxn_3_io_in_3),
    .io_out(Muxn_3_io_out)
  );
  Muxn_148 Muxn_4 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_in_3(Muxn_4_io_in_3),
    .io_out(Muxn_4_io_out)
  );
  Muxn_148 Muxn_5 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_in_3(Muxn_5_io_in_3),
    .io_out(Muxn_5_io_out)
  );
  Muxn_147 Muxn_6 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_in_4(Muxn_6_io_in_4),
    .io_out(Muxn_6_io_out)
  );
  Muxn_147 Muxn_7 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_in_4(Muxn_7_io_in_4),
    .io_out(Muxn_7_io_out)
  );
  Muxn_147 Muxn_8 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_147 Muxn_9 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNE_0 = Muxn_2_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinNE_1 = Muxn_3_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinSE_0 = Muxn_4_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSW_0 = Muxn_5_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_otrackW_0 = Muxn_6_io_out; // @[Interconnect.scala 430:21 Interconnect.scala 479:45]
  assign io_otrackN_0 = Muxn_7_io_out; // @[Interconnect.scala 431:21 Interconnect.scala 479:45]
  assign io_otrackE_0 = Muxn_8_io_out; // @[Interconnect.scala 432:21 Interconnect.scala 479:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 464:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 466:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 483:23]
  assign Muxn_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_3 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 483:23]
  assign Muxn_1_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_3 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 483:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_3 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 483:23]
  assign Muxn_3_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_3 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 483:23]
  assign Muxn_4_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 483:23]
  assign Muxn_5_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[14:12]; // @[Interconnect.scala 483:23]
  assign Muxn_6_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_4 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[17:15]; // @[Interconnect.scala 483:23]
  assign Muxn_7_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_4 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[20:18]; // @[Interconnect.scala 483:23]
  assign Muxn_8_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_4 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[23:21]; // @[Interconnect.scala 483:23]
  assign Muxn_9_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_4 = io_itrackE_0; // @[Interconnect.scala 475:63]
endmodule
module GIB_77(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire  ConfigMem_clock; // @[Interconnect.scala 463:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 463:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 463:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 463:21]
  wire [23:0] ConfigMem_io_out_0; // @[Interconnect.scala 463:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_6_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_7_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 473:25]
  wire  _T_1 = 10'ha8 == io_cfg_addr[11:2]; // @[Interconnect.scala 464:50]
  reg [31:0] _T_10; // @[Interconnect.scala 477:55]
  reg [31:0] _T_12; // @[Interconnect.scala 477:55]
  reg [31:0] _T_14; // @[Interconnect.scala 477:55]
  ConfigMem_81 ConfigMem ( // @[Interconnect.scala 463:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_148 Muxn ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_out(Muxn_io_out)
  );
  Muxn_148 Muxn_1 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_out(Muxn_1_io_out)
  );
  Muxn_148 Muxn_2 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_in_3(Muxn_2_io_in_3),
    .io_out(Muxn_2_io_out)
  );
  Muxn_148 Muxn_3 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_in_3(Muxn_3_io_in_3),
    .io_out(Muxn_3_io_out)
  );
  Muxn_148 Muxn_4 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_in_3(Muxn_4_io_in_3),
    .io_out(Muxn_4_io_out)
  );
  Muxn_148 Muxn_5 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_in_3(Muxn_5_io_in_3),
    .io_out(Muxn_5_io_out)
  );
  Muxn_147 Muxn_6 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_in_4(Muxn_6_io_in_4),
    .io_out(Muxn_6_io_out)
  );
  Muxn_147 Muxn_7 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_in_4(Muxn_7_io_in_4),
    .io_out(Muxn_7_io_out)
  );
  Muxn_147 Muxn_8 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_147 Muxn_9 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNE_0 = Muxn_2_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinNE_1 = Muxn_3_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinSE_0 = Muxn_4_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSW_0 = Muxn_5_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_otrackW_0 = _T_10; // @[Interconnect.scala 430:21 Interconnect.scala 477:45]
  assign io_otrackN_0 = _T_12; // @[Interconnect.scala 431:21 Interconnect.scala 477:45]
  assign io_otrackE_0 = _T_14; // @[Interconnect.scala 432:21 Interconnect.scala 477:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 464:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 466:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 483:23]
  assign Muxn_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_3 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 483:23]
  assign Muxn_1_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_3 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 483:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_3 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 483:23]
  assign Muxn_3_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_3 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 483:23]
  assign Muxn_4_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 483:23]
  assign Muxn_5_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[14:12]; // @[Interconnect.scala 483:23]
  assign Muxn_6_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_4 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[17:15]; // @[Interconnect.scala 483:23]
  assign Muxn_7_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_4 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[20:18]; // @[Interconnect.scala 483:23]
  assign Muxn_8_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_4 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[23:21]; // @[Interconnect.scala 483:23]
  assign Muxn_9_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_4 = io_itrackE_0; // @[Interconnect.scala 475:63]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_10 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  _T_12 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  _T_14 = _RAND_2[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_10 <= Muxn_6_io_out;
    _T_12 <= Muxn_7_io_out;
    _T_14 <= Muxn_8_io_out;
  end
endmodule
module GIB_78(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0
);
  wire  ConfigMem_clock; // @[Interconnect.scala 463:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 463:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 463:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 463:21]
  wire [23:0] ConfigMem_io_out_0; // @[Interconnect.scala 463:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_6_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_7_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 473:25]
  wire  _T_1 = 10'ha9 == io_cfg_addr[11:2]; // @[Interconnect.scala 464:50]
  ConfigMem_81 ConfigMem ( // @[Interconnect.scala 463:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_148 Muxn ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_out(Muxn_io_out)
  );
  Muxn_148 Muxn_1 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_out(Muxn_1_io_out)
  );
  Muxn_148 Muxn_2 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_in_3(Muxn_2_io_in_3),
    .io_out(Muxn_2_io_out)
  );
  Muxn_148 Muxn_3 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_in_3(Muxn_3_io_in_3),
    .io_out(Muxn_3_io_out)
  );
  Muxn_148 Muxn_4 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_in_3(Muxn_4_io_in_3),
    .io_out(Muxn_4_io_out)
  );
  Muxn_148 Muxn_5 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_in_3(Muxn_5_io_in_3),
    .io_out(Muxn_5_io_out)
  );
  Muxn_147 Muxn_6 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_in_4(Muxn_6_io_in_4),
    .io_out(Muxn_6_io_out)
  );
  Muxn_147 Muxn_7 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_in_4(Muxn_7_io_in_4),
    .io_out(Muxn_7_io_out)
  );
  Muxn_147 Muxn_8 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_147 Muxn_9 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNE_0 = Muxn_2_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinNE_1 = Muxn_3_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinSE_0 = Muxn_4_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSW_0 = Muxn_5_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_otrackW_0 = Muxn_6_io_out; // @[Interconnect.scala 430:21 Interconnect.scala 479:45]
  assign io_otrackN_0 = Muxn_7_io_out; // @[Interconnect.scala 431:21 Interconnect.scala 479:45]
  assign io_otrackE_0 = Muxn_8_io_out; // @[Interconnect.scala 432:21 Interconnect.scala 479:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 464:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 466:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 483:23]
  assign Muxn_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_3 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 483:23]
  assign Muxn_1_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_3 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 483:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_3 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 483:23]
  assign Muxn_3_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_3 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 483:23]
  assign Muxn_4_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 483:23]
  assign Muxn_5_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[14:12]; // @[Interconnect.scala 483:23]
  assign Muxn_6_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_4 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[17:15]; // @[Interconnect.scala 483:23]
  assign Muxn_7_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_4 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[20:18]; // @[Interconnect.scala 483:23]
  assign Muxn_8_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_4 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[23:21]; // @[Interconnect.scala 483:23]
  assign Muxn_9_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_4 = io_itrackE_0; // @[Interconnect.scala 475:63]
endmodule
module GIB_79(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire  ConfigMem_clock; // @[Interconnect.scala 463:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 463:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 463:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 463:21]
  wire [23:0] ConfigMem_io_out_0; // @[Interconnect.scala 463:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_6_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_7_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 473:25]
  wire  _T_1 = 10'haa == io_cfg_addr[11:2]; // @[Interconnect.scala 464:50]
  reg [31:0] _T_10; // @[Interconnect.scala 477:55]
  reg [31:0] _T_12; // @[Interconnect.scala 477:55]
  reg [31:0] _T_14; // @[Interconnect.scala 477:55]
  ConfigMem_81 ConfigMem ( // @[Interconnect.scala 463:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_148 Muxn ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_out(Muxn_io_out)
  );
  Muxn_148 Muxn_1 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_out(Muxn_1_io_out)
  );
  Muxn_148 Muxn_2 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_in_3(Muxn_2_io_in_3),
    .io_out(Muxn_2_io_out)
  );
  Muxn_148 Muxn_3 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_in_3(Muxn_3_io_in_3),
    .io_out(Muxn_3_io_out)
  );
  Muxn_148 Muxn_4 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_in_3(Muxn_4_io_in_3),
    .io_out(Muxn_4_io_out)
  );
  Muxn_148 Muxn_5 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_in_3(Muxn_5_io_in_3),
    .io_out(Muxn_5_io_out)
  );
  Muxn_147 Muxn_6 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_in_4(Muxn_6_io_in_4),
    .io_out(Muxn_6_io_out)
  );
  Muxn_147 Muxn_7 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_in_4(Muxn_7_io_in_4),
    .io_out(Muxn_7_io_out)
  );
  Muxn_147 Muxn_8 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_147 Muxn_9 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNE_0 = Muxn_2_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinNE_1 = Muxn_3_io_out; // @[Interconnect.scala 427:20 Interconnect.scala 479:45]
  assign io_ipinSE_0 = Muxn_4_io_out; // @[Interconnect.scala 429:20 Interconnect.scala 479:45]
  assign io_ipinSW_0 = Muxn_5_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_otrackW_0 = _T_10; // @[Interconnect.scala 430:21 Interconnect.scala 477:45]
  assign io_otrackN_0 = _T_12; // @[Interconnect.scala 431:21 Interconnect.scala 477:45]
  assign io_otrackE_0 = _T_14; // @[Interconnect.scala 432:21 Interconnect.scala 477:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 464:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 466:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 483:23]
  assign Muxn_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_3 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 483:23]
  assign Muxn_1_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_2 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_3 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 483:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_3 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 483:23]
  assign Muxn_3_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_3 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 483:23]
  assign Muxn_4_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 483:23]
  assign Muxn_5_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[14:12]; // @[Interconnect.scala 483:23]
  assign Muxn_6_io_in_0 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_1 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_4 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[17:15]; // @[Interconnect.scala 483:23]
  assign Muxn_7_io_in_0 = io_opinSE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_3 = io_itrackE_0; // @[Interconnect.scala 475:63]
  assign Muxn_7_io_in_4 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[20:18]; // @[Interconnect.scala 483:23]
  assign Muxn_8_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_8_io_in_4 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[23:21]; // @[Interconnect.scala 483:23]
  assign Muxn_9_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_1 = io_opinNE_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_9_io_in_4 = io_itrackE_0; // @[Interconnect.scala 475:63]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_10 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  _T_12 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  _T_14 = _RAND_2[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_10 <= Muxn_6_io_out;
    _T_12 <= Muxn_7_io_out;
    _T_14 <= Muxn_8_io_out;
  end
endmodule
module GIB_80(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinSW_0,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0
);
  wire  ConfigMem_clock; // @[Interconnect.scala 463:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 463:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 463:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 463:21]
  wire [13:0] ConfigMem_io_out_0; // @[Interconnect.scala 463:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 473:25]
  wire  Muxn_2_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 473:25]
  wire [2:0] Muxn_5_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_in_4; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 473:25]
  wire [1:0] Muxn_6_io_config; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 473:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 473:25]
  wire  _T_1 = 10'hab == io_cfg_addr[11:2]; // @[Interconnect.scala 464:50]
  ConfigMem_80 ConfigMem ( // @[Interconnect.scala 463:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_145 Muxn ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_out(Muxn_io_out)
  );
  Muxn_145 Muxn_1 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_out(Muxn_1_io_out)
  );
  Muxn Muxn_2 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_out(Muxn_2_io_out)
  );
  Muxn_145 Muxn_3 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_out(Muxn_3_io_out)
  );
  Muxn_148 Muxn_4 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_in_3(Muxn_4_io_in_3),
    .io_out(Muxn_4_io_out)
  );
  Muxn_147 Muxn_5 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_in_3(Muxn_5_io_in_3),
    .io_in_4(Muxn_5_io_in_4),
    .io_out(Muxn_5_io_out)
  );
  Muxn_148 Muxn_6 ( // @[Interconnect.scala 473:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_out(Muxn_6_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 426:20 Interconnect.scala 479:45]
  assign io_ipinSW_0 = Muxn_2_io_out; // @[Interconnect.scala 428:20 Interconnect.scala 479:45]
  assign io_otrackW_0 = Muxn_3_io_out; // @[Interconnect.scala 430:21 Interconnect.scala 479:45]
  assign io_otrackN_0 = Muxn_4_io_out; // @[Interconnect.scala 431:21 Interconnect.scala 479:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 464:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 466:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 483:23]
  assign Muxn_io_in_0 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_1 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_io_in_2 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 483:23]
  assign Muxn_1_io_in_0 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_1 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_1_io_in_2 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[4]; // @[Interconnect.scala 483:23]
  assign Muxn_2_io_in_0 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_2_io_in_1 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[6:5]; // @[Interconnect.scala 483:23]
  assign Muxn_3_io_in_0 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_1 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_3_io_in_2 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[8:7]; // @[Interconnect.scala 483:23]
  assign Muxn_4_io_in_0 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_1 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_2 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_4_io_in_3 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:9]; // @[Interconnect.scala 483:23]
  assign Muxn_5_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_1 = io_opinSW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_2 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_3 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_5_io_in_4 = 32'h0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[13:12]; // @[Interconnect.scala 483:23]
  assign Muxn_6_io_in_0 = io_opinNW_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_1 = io_itrackW_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_2 = io_itrackN_0; // @[Interconnect.scala 475:63]
  assign Muxn_6_io_in_3 = 32'h0; // @[Interconnect.scala 475:63]
endmodule
module CGRA(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [11:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en_0,
  input         io_en_1,
  input         io_en_2,
  input         io_en_3,
  input         io_en_4,
  input         io_en_5,
  input         io_en_6,
  input         io_en_7,
  input         io_en_8,
  input         io_en_9,
  input         io_en_10,
  input         io_en_11,
  input         io_en_12,
  input         io_en_13,
  input         io_en_14,
  input         io_en_15,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  input  [31:0] io_in_8,
  input  [31:0] io_in_9,
  input  [31:0] io_in_10,
  input  [31:0] io_in_11,
  input  [31:0] io_in_12,
  input  [31:0] io_in_13,
  input  [31:0] io_in_14,
  input  [31:0] io_in_15,
  output [31:0] io_out_0,
  output [31:0] io_out_1,
  output [31:0] io_out_2,
  output [31:0] io_out_3,
  output [31:0] io_out_4,
  output [31:0] io_out_5,
  output [31:0] io_out_6,
  output [31:0] io_out_7,
  output [31:0] io_out_8,
  output [31:0] io_out_9,
  output [31:0] io_out_10,
  output [31:0] io_out_11,
  output [31:0] io_out_12,
  output [31:0] io_out_13,
  output [31:0] io_out_14,
  output [31:0] io_out_15
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_19;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] ibs_0_io_in_0; // @[CGRA.scala 149:20]
  wire [31:0] ibs_0_io_out_0; // @[CGRA.scala 149:20]
  wire [31:0] ibs_1_io_in_0; // @[CGRA.scala 149:20]
  wire [31:0] ibs_1_io_out_0; // @[CGRA.scala 149:20]
  wire [31:0] ibs_2_io_in_0; // @[CGRA.scala 149:20]
  wire [31:0] ibs_2_io_out_0; // @[CGRA.scala 149:20]
  wire [31:0] ibs_3_io_in_0; // @[CGRA.scala 149:20]
  wire [31:0] ibs_3_io_out_0; // @[CGRA.scala 149:20]
  wire [31:0] ibs_4_io_in_0; // @[CGRA.scala 149:20]
  wire [31:0] ibs_4_io_out_0; // @[CGRA.scala 149:20]
  wire [31:0] ibs_5_io_in_0; // @[CGRA.scala 149:20]
  wire [31:0] ibs_5_io_out_0; // @[CGRA.scala 149:20]
  wire [31:0] ibs_6_io_in_0; // @[CGRA.scala 149:20]
  wire [31:0] ibs_6_io_out_0; // @[CGRA.scala 149:20]
  wire [31:0] ibs_7_io_in_0; // @[CGRA.scala 149:20]
  wire [31:0] ibs_7_io_out_0; // @[CGRA.scala 149:20]
  wire [31:0] ibs_8_io_in_0; // @[CGRA.scala 149:20]
  wire [31:0] ibs_8_io_out_0; // @[CGRA.scala 149:20]
  wire [31:0] ibs_9_io_in_0; // @[CGRA.scala 149:20]
  wire [31:0] ibs_9_io_out_0; // @[CGRA.scala 149:20]
  wire [31:0] ibs_10_io_in_0; // @[CGRA.scala 149:20]
  wire [31:0] ibs_10_io_out_0; // @[CGRA.scala 149:20]
  wire [31:0] ibs_11_io_in_0; // @[CGRA.scala 149:20]
  wire [31:0] ibs_11_io_out_0; // @[CGRA.scala 149:20]
  wire [31:0] ibs_12_io_in_0; // @[CGRA.scala 149:20]
  wire [31:0] ibs_12_io_out_0; // @[CGRA.scala 149:20]
  wire [31:0] ibs_13_io_in_0; // @[CGRA.scala 149:20]
  wire [31:0] ibs_13_io_out_0; // @[CGRA.scala 149:20]
  wire [31:0] ibs_14_io_in_0; // @[CGRA.scala 149:20]
  wire [31:0] ibs_14_io_out_0; // @[CGRA.scala 149:20]
  wire [31:0] ibs_15_io_in_0; // @[CGRA.scala 149:20]
  wire [31:0] ibs_15_io_out_0; // @[CGRA.scala 149:20]
  wire  obs_0_clock; // @[CGRA.scala 176:20]
  wire  obs_0_reset; // @[CGRA.scala 176:20]
  wire  obs_0_io_cfg_en; // @[CGRA.scala 176:20]
  wire [11:0] obs_0_io_cfg_addr; // @[CGRA.scala 176:20]
  wire [31:0] obs_0_io_cfg_data; // @[CGRA.scala 176:20]
  wire [31:0] obs_0_io_in_0; // @[CGRA.scala 176:20]
  wire [31:0] obs_0_io_in_1; // @[CGRA.scala 176:20]
  wire [31:0] obs_0_io_out_0; // @[CGRA.scala 176:20]
  wire  obs_1_clock; // @[CGRA.scala 176:20]
  wire  obs_1_reset; // @[CGRA.scala 176:20]
  wire  obs_1_io_cfg_en; // @[CGRA.scala 176:20]
  wire [11:0] obs_1_io_cfg_addr; // @[CGRA.scala 176:20]
  wire [31:0] obs_1_io_cfg_data; // @[CGRA.scala 176:20]
  wire [31:0] obs_1_io_in_0; // @[CGRA.scala 176:20]
  wire [31:0] obs_1_io_in_1; // @[CGRA.scala 176:20]
  wire [31:0] obs_1_io_out_0; // @[CGRA.scala 176:20]
  wire  obs_2_clock; // @[CGRA.scala 176:20]
  wire  obs_2_reset; // @[CGRA.scala 176:20]
  wire  obs_2_io_cfg_en; // @[CGRA.scala 176:20]
  wire [11:0] obs_2_io_cfg_addr; // @[CGRA.scala 176:20]
  wire [31:0] obs_2_io_cfg_data; // @[CGRA.scala 176:20]
  wire [31:0] obs_2_io_in_0; // @[CGRA.scala 176:20]
  wire [31:0] obs_2_io_in_1; // @[CGRA.scala 176:20]
  wire [31:0] obs_2_io_out_0; // @[CGRA.scala 176:20]
  wire  obs_3_clock; // @[CGRA.scala 176:20]
  wire  obs_3_reset; // @[CGRA.scala 176:20]
  wire  obs_3_io_cfg_en; // @[CGRA.scala 176:20]
  wire [11:0] obs_3_io_cfg_addr; // @[CGRA.scala 176:20]
  wire [31:0] obs_3_io_cfg_data; // @[CGRA.scala 176:20]
  wire [31:0] obs_3_io_in_0; // @[CGRA.scala 176:20]
  wire [31:0] obs_3_io_in_1; // @[CGRA.scala 176:20]
  wire [31:0] obs_3_io_out_0; // @[CGRA.scala 176:20]
  wire  obs_4_clock; // @[CGRA.scala 176:20]
  wire  obs_4_reset; // @[CGRA.scala 176:20]
  wire  obs_4_io_cfg_en; // @[CGRA.scala 176:20]
  wire [11:0] obs_4_io_cfg_addr; // @[CGRA.scala 176:20]
  wire [31:0] obs_4_io_cfg_data; // @[CGRA.scala 176:20]
  wire [31:0] obs_4_io_in_0; // @[CGRA.scala 176:20]
  wire [31:0] obs_4_io_in_1; // @[CGRA.scala 176:20]
  wire [31:0] obs_4_io_out_0; // @[CGRA.scala 176:20]
  wire  obs_5_clock; // @[CGRA.scala 176:20]
  wire  obs_5_reset; // @[CGRA.scala 176:20]
  wire  obs_5_io_cfg_en; // @[CGRA.scala 176:20]
  wire [11:0] obs_5_io_cfg_addr; // @[CGRA.scala 176:20]
  wire [31:0] obs_5_io_cfg_data; // @[CGRA.scala 176:20]
  wire [31:0] obs_5_io_in_0; // @[CGRA.scala 176:20]
  wire [31:0] obs_5_io_in_1; // @[CGRA.scala 176:20]
  wire [31:0] obs_5_io_out_0; // @[CGRA.scala 176:20]
  wire  obs_6_clock; // @[CGRA.scala 176:20]
  wire  obs_6_reset; // @[CGRA.scala 176:20]
  wire  obs_6_io_cfg_en; // @[CGRA.scala 176:20]
  wire [11:0] obs_6_io_cfg_addr; // @[CGRA.scala 176:20]
  wire [31:0] obs_6_io_cfg_data; // @[CGRA.scala 176:20]
  wire [31:0] obs_6_io_in_0; // @[CGRA.scala 176:20]
  wire [31:0] obs_6_io_in_1; // @[CGRA.scala 176:20]
  wire [31:0] obs_6_io_out_0; // @[CGRA.scala 176:20]
  wire  obs_7_clock; // @[CGRA.scala 176:20]
  wire  obs_7_reset; // @[CGRA.scala 176:20]
  wire  obs_7_io_cfg_en; // @[CGRA.scala 176:20]
  wire [11:0] obs_7_io_cfg_addr; // @[CGRA.scala 176:20]
  wire [31:0] obs_7_io_cfg_data; // @[CGRA.scala 176:20]
  wire [31:0] obs_7_io_in_0; // @[CGRA.scala 176:20]
  wire [31:0] obs_7_io_in_1; // @[CGRA.scala 176:20]
  wire [31:0] obs_7_io_out_0; // @[CGRA.scala 176:20]
  wire  obs_8_clock; // @[CGRA.scala 176:20]
  wire  obs_8_reset; // @[CGRA.scala 176:20]
  wire  obs_8_io_cfg_en; // @[CGRA.scala 176:20]
  wire [11:0] obs_8_io_cfg_addr; // @[CGRA.scala 176:20]
  wire [31:0] obs_8_io_cfg_data; // @[CGRA.scala 176:20]
  wire [31:0] obs_8_io_in_0; // @[CGRA.scala 176:20]
  wire [31:0] obs_8_io_in_1; // @[CGRA.scala 176:20]
  wire [31:0] obs_8_io_out_0; // @[CGRA.scala 176:20]
  wire  obs_9_clock; // @[CGRA.scala 176:20]
  wire  obs_9_reset; // @[CGRA.scala 176:20]
  wire  obs_9_io_cfg_en; // @[CGRA.scala 176:20]
  wire [11:0] obs_9_io_cfg_addr; // @[CGRA.scala 176:20]
  wire [31:0] obs_9_io_cfg_data; // @[CGRA.scala 176:20]
  wire [31:0] obs_9_io_in_0; // @[CGRA.scala 176:20]
  wire [31:0] obs_9_io_in_1; // @[CGRA.scala 176:20]
  wire [31:0] obs_9_io_out_0; // @[CGRA.scala 176:20]
  wire  obs_10_clock; // @[CGRA.scala 176:20]
  wire  obs_10_reset; // @[CGRA.scala 176:20]
  wire  obs_10_io_cfg_en; // @[CGRA.scala 176:20]
  wire [11:0] obs_10_io_cfg_addr; // @[CGRA.scala 176:20]
  wire [31:0] obs_10_io_cfg_data; // @[CGRA.scala 176:20]
  wire [31:0] obs_10_io_in_0; // @[CGRA.scala 176:20]
  wire [31:0] obs_10_io_in_1; // @[CGRA.scala 176:20]
  wire [31:0] obs_10_io_out_0; // @[CGRA.scala 176:20]
  wire  obs_11_clock; // @[CGRA.scala 176:20]
  wire  obs_11_reset; // @[CGRA.scala 176:20]
  wire  obs_11_io_cfg_en; // @[CGRA.scala 176:20]
  wire [11:0] obs_11_io_cfg_addr; // @[CGRA.scala 176:20]
  wire [31:0] obs_11_io_cfg_data; // @[CGRA.scala 176:20]
  wire [31:0] obs_11_io_in_0; // @[CGRA.scala 176:20]
  wire [31:0] obs_11_io_in_1; // @[CGRA.scala 176:20]
  wire [31:0] obs_11_io_out_0; // @[CGRA.scala 176:20]
  wire  obs_12_clock; // @[CGRA.scala 176:20]
  wire  obs_12_reset; // @[CGRA.scala 176:20]
  wire  obs_12_io_cfg_en; // @[CGRA.scala 176:20]
  wire [11:0] obs_12_io_cfg_addr; // @[CGRA.scala 176:20]
  wire [31:0] obs_12_io_cfg_data; // @[CGRA.scala 176:20]
  wire [31:0] obs_12_io_in_0; // @[CGRA.scala 176:20]
  wire [31:0] obs_12_io_in_1; // @[CGRA.scala 176:20]
  wire [31:0] obs_12_io_out_0; // @[CGRA.scala 176:20]
  wire  obs_13_clock; // @[CGRA.scala 176:20]
  wire  obs_13_reset; // @[CGRA.scala 176:20]
  wire  obs_13_io_cfg_en; // @[CGRA.scala 176:20]
  wire [11:0] obs_13_io_cfg_addr; // @[CGRA.scala 176:20]
  wire [31:0] obs_13_io_cfg_data; // @[CGRA.scala 176:20]
  wire [31:0] obs_13_io_in_0; // @[CGRA.scala 176:20]
  wire [31:0] obs_13_io_in_1; // @[CGRA.scala 176:20]
  wire [31:0] obs_13_io_out_0; // @[CGRA.scala 176:20]
  wire  obs_14_clock; // @[CGRA.scala 176:20]
  wire  obs_14_reset; // @[CGRA.scala 176:20]
  wire  obs_14_io_cfg_en; // @[CGRA.scala 176:20]
  wire [11:0] obs_14_io_cfg_addr; // @[CGRA.scala 176:20]
  wire [31:0] obs_14_io_cfg_data; // @[CGRA.scala 176:20]
  wire [31:0] obs_14_io_in_0; // @[CGRA.scala 176:20]
  wire [31:0] obs_14_io_in_1; // @[CGRA.scala 176:20]
  wire [31:0] obs_14_io_out_0; // @[CGRA.scala 176:20]
  wire  obs_15_clock; // @[CGRA.scala 176:20]
  wire  obs_15_reset; // @[CGRA.scala 176:20]
  wire  obs_15_io_cfg_en; // @[CGRA.scala 176:20]
  wire [11:0] obs_15_io_cfg_addr; // @[CGRA.scala 176:20]
  wire [31:0] obs_15_io_cfg_data; // @[CGRA.scala 176:20]
  wire [31:0] obs_15_io_in_0; // @[CGRA.scala 176:20]
  wire [31:0] obs_15_io_in_1; // @[CGRA.scala 176:20]
  wire [31:0] obs_15_io_out_0; // @[CGRA.scala 176:20]
  wire  pes_0_clock; // @[CGRA.scala 200:20]
  wire  pes_0_reset; // @[CGRA.scala 200:20]
  wire  pes_0_io_cfg_en; // @[CGRA.scala 200:20]
  wire [11:0] pes_0_io_cfg_addr; // @[CGRA.scala 200:20]
  wire [31:0] pes_0_io_cfg_data; // @[CGRA.scala 200:20]
  wire  pes_0_io_en; // @[CGRA.scala 200:20]
  wire [31:0] pes_0_io_in_0; // @[CGRA.scala 200:20]
  wire [31:0] pes_0_io_in_1; // @[CGRA.scala 200:20]
  wire [31:0] pes_0_io_in_2; // @[CGRA.scala 200:20]
  wire [31:0] pes_0_io_in_3; // @[CGRA.scala 200:20]
  wire [31:0] pes_0_io_in_4; // @[CGRA.scala 200:20]
  wire [31:0] pes_0_io_in_5; // @[CGRA.scala 200:20]
  wire [31:0] pes_0_io_in_6; // @[CGRA.scala 200:20]
  wire [31:0] pes_0_io_in_7; // @[CGRA.scala 200:20]
  wire [31:0] pes_0_io_out_0; // @[CGRA.scala 200:20]
  wire  pes_1_clock; // @[CGRA.scala 200:20]
  wire  pes_1_reset; // @[CGRA.scala 200:20]
  wire  pes_1_io_cfg_en; // @[CGRA.scala 200:20]
  wire [11:0] pes_1_io_cfg_addr; // @[CGRA.scala 200:20]
  wire [31:0] pes_1_io_cfg_data; // @[CGRA.scala 200:20]
  wire  pes_1_io_en; // @[CGRA.scala 200:20]
  wire [31:0] pes_1_io_in_0; // @[CGRA.scala 200:20]
  wire [31:0] pes_1_io_in_1; // @[CGRA.scala 200:20]
  wire [31:0] pes_1_io_in_2; // @[CGRA.scala 200:20]
  wire [31:0] pes_1_io_in_3; // @[CGRA.scala 200:20]
  wire [31:0] pes_1_io_in_4; // @[CGRA.scala 200:20]
  wire [31:0] pes_1_io_in_5; // @[CGRA.scala 200:20]
  wire [31:0] pes_1_io_in_6; // @[CGRA.scala 200:20]
  wire [31:0] pes_1_io_in_7; // @[CGRA.scala 200:20]
  wire [31:0] pes_1_io_out_0; // @[CGRA.scala 200:20]
  wire  pes_2_clock; // @[CGRA.scala 200:20]
  wire  pes_2_reset; // @[CGRA.scala 200:20]
  wire  pes_2_io_cfg_en; // @[CGRA.scala 200:20]
  wire [11:0] pes_2_io_cfg_addr; // @[CGRA.scala 200:20]
  wire [31:0] pes_2_io_cfg_data; // @[CGRA.scala 200:20]
  wire  pes_2_io_en; // @[CGRA.scala 200:20]
  wire [31:0] pes_2_io_in_0; // @[CGRA.scala 200:20]
  wire [31:0] pes_2_io_in_1; // @[CGRA.scala 200:20]
  wire [31:0] pes_2_io_in_2; // @[CGRA.scala 200:20]
  wire [31:0] pes_2_io_in_3; // @[CGRA.scala 200:20]
  wire [31:0] pes_2_io_in_4; // @[CGRA.scala 200:20]
  wire [31:0] pes_2_io_in_5; // @[CGRA.scala 200:20]
  wire [31:0] pes_2_io_in_6; // @[CGRA.scala 200:20]
  wire [31:0] pes_2_io_in_7; // @[CGRA.scala 200:20]
  wire [31:0] pes_2_io_out_0; // @[CGRA.scala 200:20]
  wire  pes_3_clock; // @[CGRA.scala 200:20]
  wire  pes_3_reset; // @[CGRA.scala 200:20]
  wire  pes_3_io_cfg_en; // @[CGRA.scala 200:20]
  wire [11:0] pes_3_io_cfg_addr; // @[CGRA.scala 200:20]
  wire [31:0] pes_3_io_cfg_data; // @[CGRA.scala 200:20]
  wire  pes_3_io_en; // @[CGRA.scala 200:20]
  wire [31:0] pes_3_io_in_0; // @[CGRA.scala 200:20]
  wire [31:0] pes_3_io_in_1; // @[CGRA.scala 200:20]
  wire [31:0] pes_3_io_in_2; // @[CGRA.scala 200:20]
  wire [31:0] pes_3_io_in_3; // @[CGRA.scala 200:20]
  wire [31:0] pes_3_io_in_4; // @[CGRA.scala 200:20]
  wire [31:0] pes_3_io_in_5; // @[CGRA.scala 200:20]
  wire [31:0] pes_3_io_in_6; // @[CGRA.scala 200:20]
  wire [31:0] pes_3_io_in_7; // @[CGRA.scala 200:20]
  wire [31:0] pes_3_io_out_0; // @[CGRA.scala 200:20]
  wire  pes_4_clock; // @[CGRA.scala 200:20]
  wire  pes_4_reset; // @[CGRA.scala 200:20]
  wire  pes_4_io_cfg_en; // @[CGRA.scala 200:20]
  wire [11:0] pes_4_io_cfg_addr; // @[CGRA.scala 200:20]
  wire [31:0] pes_4_io_cfg_data; // @[CGRA.scala 200:20]
  wire  pes_4_io_en; // @[CGRA.scala 200:20]
  wire [31:0] pes_4_io_in_0; // @[CGRA.scala 200:20]
  wire [31:0] pes_4_io_in_1; // @[CGRA.scala 200:20]
  wire [31:0] pes_4_io_in_2; // @[CGRA.scala 200:20]
  wire [31:0] pes_4_io_in_3; // @[CGRA.scala 200:20]
  wire [31:0] pes_4_io_in_4; // @[CGRA.scala 200:20]
  wire [31:0] pes_4_io_in_5; // @[CGRA.scala 200:20]
  wire [31:0] pes_4_io_in_6; // @[CGRA.scala 200:20]
  wire [31:0] pes_4_io_in_7; // @[CGRA.scala 200:20]
  wire [31:0] pes_4_io_out_0; // @[CGRA.scala 200:20]
  wire  pes_5_clock; // @[CGRA.scala 200:20]
  wire  pes_5_reset; // @[CGRA.scala 200:20]
  wire  pes_5_io_cfg_en; // @[CGRA.scala 200:20]
  wire [11:0] pes_5_io_cfg_addr; // @[CGRA.scala 200:20]
  wire [31:0] pes_5_io_cfg_data; // @[CGRA.scala 200:20]
  wire  pes_5_io_en; // @[CGRA.scala 200:20]
  wire [31:0] pes_5_io_in_0; // @[CGRA.scala 200:20]
  wire [31:0] pes_5_io_in_1; // @[CGRA.scala 200:20]
  wire [31:0] pes_5_io_in_2; // @[CGRA.scala 200:20]
  wire [31:0] pes_5_io_in_3; // @[CGRA.scala 200:20]
  wire [31:0] pes_5_io_in_4; // @[CGRA.scala 200:20]
  wire [31:0] pes_5_io_in_5; // @[CGRA.scala 200:20]
  wire [31:0] pes_5_io_in_6; // @[CGRA.scala 200:20]
  wire [31:0] pes_5_io_in_7; // @[CGRA.scala 200:20]
  wire [31:0] pes_5_io_out_0; // @[CGRA.scala 200:20]
  wire  pes_6_clock; // @[CGRA.scala 200:20]
  wire  pes_6_reset; // @[CGRA.scala 200:20]
  wire  pes_6_io_cfg_en; // @[CGRA.scala 200:20]
  wire [11:0] pes_6_io_cfg_addr; // @[CGRA.scala 200:20]
  wire [31:0] pes_6_io_cfg_data; // @[CGRA.scala 200:20]
  wire  pes_6_io_en; // @[CGRA.scala 200:20]
  wire [31:0] pes_6_io_in_0; // @[CGRA.scala 200:20]
  wire [31:0] pes_6_io_in_1; // @[CGRA.scala 200:20]
  wire [31:0] pes_6_io_in_2; // @[CGRA.scala 200:20]
  wire [31:0] pes_6_io_in_3; // @[CGRA.scala 200:20]
  wire [31:0] pes_6_io_in_4; // @[CGRA.scala 200:20]
  wire [31:0] pes_6_io_in_5; // @[CGRA.scala 200:20]
  wire [31:0] pes_6_io_in_6; // @[CGRA.scala 200:20]
  wire [31:0] pes_6_io_in_7; // @[CGRA.scala 200:20]
  wire [31:0] pes_6_io_out_0; // @[CGRA.scala 200:20]
  wire  pes_7_clock; // @[CGRA.scala 200:20]
  wire  pes_7_reset; // @[CGRA.scala 200:20]
  wire  pes_7_io_cfg_en; // @[CGRA.scala 200:20]
  wire [11:0] pes_7_io_cfg_addr; // @[CGRA.scala 200:20]
  wire [31:0] pes_7_io_cfg_data; // @[CGRA.scala 200:20]
  wire  pes_7_io_en; // @[CGRA.scala 200:20]
  wire [31:0] pes_7_io_in_0; // @[CGRA.scala 200:20]
  wire [31:0] pes_7_io_in_1; // @[CGRA.scala 200:20]
  wire [31:0] pes_7_io_in_2; // @[CGRA.scala 200:20]
  wire [31:0] pes_7_io_in_3; // @[CGRA.scala 200:20]
  wire [31:0] pes_7_io_in_4; // @[CGRA.scala 200:20]
  wire [31:0] pes_7_io_in_5; // @[CGRA.scala 200:20]
  wire [31:0] pes_7_io_in_6; // @[CGRA.scala 200:20]
  wire [31:0] pes_7_io_in_7; // @[CGRA.scala 200:20]
  wire [31:0] pes_7_io_out_0; // @[CGRA.scala 200:20]
  wire  pes_8_clock; // @[CGRA.scala 200:20]
  wire  pes_8_reset; // @[CGRA.scala 200:20]
  wire  pes_8_io_cfg_en; // @[CGRA.scala 200:20]
  wire [11:0] pes_8_io_cfg_addr; // @[CGRA.scala 200:20]
  wire [31:0] pes_8_io_cfg_data; // @[CGRA.scala 200:20]
  wire  pes_8_io_en; // @[CGRA.scala 200:20]
  wire [31:0] pes_8_io_in_0; // @[CGRA.scala 200:20]
  wire [31:0] pes_8_io_in_1; // @[CGRA.scala 200:20]
  wire [31:0] pes_8_io_in_2; // @[CGRA.scala 200:20]
  wire [31:0] pes_8_io_in_3; // @[CGRA.scala 200:20]
  wire [31:0] pes_8_io_in_4; // @[CGRA.scala 200:20]
  wire [31:0] pes_8_io_in_5; // @[CGRA.scala 200:20]
  wire [31:0] pes_8_io_in_6; // @[CGRA.scala 200:20]
  wire [31:0] pes_8_io_in_7; // @[CGRA.scala 200:20]
  wire [31:0] pes_8_io_out_0; // @[CGRA.scala 200:20]
  wire  pes_9_clock; // @[CGRA.scala 200:20]
  wire  pes_9_reset; // @[CGRA.scala 200:20]
  wire  pes_9_io_cfg_en; // @[CGRA.scala 200:20]
  wire [11:0] pes_9_io_cfg_addr; // @[CGRA.scala 200:20]
  wire [31:0] pes_9_io_cfg_data; // @[CGRA.scala 200:20]
  wire  pes_9_io_en; // @[CGRA.scala 200:20]
  wire [31:0] pes_9_io_in_0; // @[CGRA.scala 200:20]
  wire [31:0] pes_9_io_in_1; // @[CGRA.scala 200:20]
  wire [31:0] pes_9_io_in_2; // @[CGRA.scala 200:20]
  wire [31:0] pes_9_io_in_3; // @[CGRA.scala 200:20]
  wire [31:0] pes_9_io_in_4; // @[CGRA.scala 200:20]
  wire [31:0] pes_9_io_in_5; // @[CGRA.scala 200:20]
  wire [31:0] pes_9_io_in_6; // @[CGRA.scala 200:20]
  wire [31:0] pes_9_io_in_7; // @[CGRA.scala 200:20]
  wire [31:0] pes_9_io_out_0; // @[CGRA.scala 200:20]
  wire  pes_10_clock; // @[CGRA.scala 200:20]
  wire  pes_10_reset; // @[CGRA.scala 200:20]
  wire  pes_10_io_cfg_en; // @[CGRA.scala 200:20]
  wire [11:0] pes_10_io_cfg_addr; // @[CGRA.scala 200:20]
  wire [31:0] pes_10_io_cfg_data; // @[CGRA.scala 200:20]
  wire  pes_10_io_en; // @[CGRA.scala 200:20]
  wire [31:0] pes_10_io_in_0; // @[CGRA.scala 200:20]
  wire [31:0] pes_10_io_in_1; // @[CGRA.scala 200:20]
  wire [31:0] pes_10_io_in_2; // @[CGRA.scala 200:20]
  wire [31:0] pes_10_io_in_3; // @[CGRA.scala 200:20]
  wire [31:0] pes_10_io_in_4; // @[CGRA.scala 200:20]
  wire [31:0] pes_10_io_in_5; // @[CGRA.scala 200:20]
  wire [31:0] pes_10_io_in_6; // @[CGRA.scala 200:20]
  wire [31:0] pes_10_io_in_7; // @[CGRA.scala 200:20]
  wire [31:0] pes_10_io_out_0; // @[CGRA.scala 200:20]
  wire  pes_11_clock; // @[CGRA.scala 200:20]
  wire  pes_11_reset; // @[CGRA.scala 200:20]
  wire  pes_11_io_cfg_en; // @[CGRA.scala 200:20]
  wire [11:0] pes_11_io_cfg_addr; // @[CGRA.scala 200:20]
  wire [31:0] pes_11_io_cfg_data; // @[CGRA.scala 200:20]
  wire  pes_11_io_en; // @[CGRA.scala 200:20]
  wire [31:0] pes_11_io_in_0; // @[CGRA.scala 200:20]
  wire [31:0] pes_11_io_in_1; // @[CGRA.scala 200:20]
  wire [31:0] pes_11_io_in_2; // @[CGRA.scala 200:20]
  wire [31:0] pes_11_io_in_3; // @[CGRA.scala 200:20]
  wire [31:0] pes_11_io_in_4; // @[CGRA.scala 200:20]
  wire [31:0] pes_11_io_in_5; // @[CGRA.scala 200:20]
  wire [31:0] pes_11_io_in_6; // @[CGRA.scala 200:20]
  wire [31:0] pes_11_io_in_7; // @[CGRA.scala 200:20]
  wire [31:0] pes_11_io_out_0; // @[CGRA.scala 200:20]
  wire  pes_12_clock; // @[CGRA.scala 200:20]
  wire  pes_12_reset; // @[CGRA.scala 200:20]
  wire  pes_12_io_cfg_en; // @[CGRA.scala 200:20]
  wire [11:0] pes_12_io_cfg_addr; // @[CGRA.scala 200:20]
  wire [31:0] pes_12_io_cfg_data; // @[CGRA.scala 200:20]
  wire  pes_12_io_en; // @[CGRA.scala 200:20]
  wire [31:0] pes_12_io_in_0; // @[CGRA.scala 200:20]
  wire [31:0] pes_12_io_in_1; // @[CGRA.scala 200:20]
  wire [31:0] pes_12_io_in_2; // @[CGRA.scala 200:20]
  wire [31:0] pes_12_io_in_3; // @[CGRA.scala 200:20]
  wire [31:0] pes_12_io_in_4; // @[CGRA.scala 200:20]
  wire [31:0] pes_12_io_in_5; // @[CGRA.scala 200:20]
  wire [31:0] pes_12_io_in_6; // @[CGRA.scala 200:20]
  wire [31:0] pes_12_io_in_7; // @[CGRA.scala 200:20]
  wire [31:0] pes_12_io_out_0; // @[CGRA.scala 200:20]
  wire  pes_13_clock; // @[CGRA.scala 200:20]
  wire  pes_13_reset; // @[CGRA.scala 200:20]
  wire  pes_13_io_cfg_en; // @[CGRA.scala 200:20]
  wire [11:0] pes_13_io_cfg_addr; // @[CGRA.scala 200:20]
  wire [31:0] pes_13_io_cfg_data; // @[CGRA.scala 200:20]
  wire  pes_13_io_en; // @[CGRA.scala 200:20]
  wire [31:0] pes_13_io_in_0; // @[CGRA.scala 200:20]
  wire [31:0] pes_13_io_in_1; // @[CGRA.scala 200:20]
  wire [31:0] pes_13_io_in_2; // @[CGRA.scala 200:20]
  wire [31:0] pes_13_io_in_3; // @[CGRA.scala 200:20]
  wire [31:0] pes_13_io_in_4; // @[CGRA.scala 200:20]
  wire [31:0] pes_13_io_in_5; // @[CGRA.scala 200:20]
  wire [31:0] pes_13_io_in_6; // @[CGRA.scala 200:20]
  wire [31:0] pes_13_io_in_7; // @[CGRA.scala 200:20]
  wire [31:0] pes_13_io_out_0; // @[CGRA.scala 200:20]
  wire  pes_14_clock; // @[CGRA.scala 200:20]
  wire  pes_14_reset; // @[CGRA.scala 200:20]
  wire  pes_14_io_cfg_en; // @[CGRA.scala 200:20]
  wire [11:0] pes_14_io_cfg_addr; // @[CGRA.scala 200:20]
  wire [31:0] pes_14_io_cfg_data; // @[CGRA.scala 200:20]
  wire  pes_14_io_en; // @[CGRA.scala 200:20]
  wire [31:0] pes_14_io_in_0; // @[CGRA.scala 200:20]
  wire [31:0] pes_14_io_in_1; // @[CGRA.scala 200:20]
  wire [31:0] pes_14_io_in_2; // @[CGRA.scala 200:20]
  wire [31:0] pes_14_io_in_3; // @[CGRA.scala 200:20]
  wire [31:0] pes_14_io_in_4; // @[CGRA.scala 200:20]
  wire [31:0] pes_14_io_in_5; // @[CGRA.scala 200:20]
  wire [31:0] pes_14_io_in_6; // @[CGRA.scala 200:20]
  wire [31:0] pes_14_io_in_7; // @[CGRA.scala 200:20]
  wire [31:0] pes_14_io_out_0; // @[CGRA.scala 200:20]
  wire  pes_15_clock; // @[CGRA.scala 200:20]
  wire  pes_15_reset; // @[CGRA.scala 200:20]
  wire  pes_15_io_cfg_en; // @[CGRA.scala 200:20]
  wire [11:0] pes_15_io_cfg_addr; // @[CGRA.scala 200:20]
  wire [31:0] pes_15_io_cfg_data; // @[CGRA.scala 200:20]
  wire  pes_15_io_en; // @[CGRA.scala 200:20]
  wire [31:0] pes_15_io_in_0; // @[CGRA.scala 200:20]
  wire [31:0] pes_15_io_in_1; // @[CGRA.scala 200:20]
  wire [31:0] pes_15_io_in_2; // @[CGRA.scala 200:20]
  wire [31:0] pes_15_io_in_3; // @[CGRA.scala 200:20]
  wire [31:0] pes_15_io_in_4; // @[CGRA.scala 200:20]
  wire [31:0] pes_15_io_in_5; // @[CGRA.scala 200:20]
  wire [31:0] pes_15_io_in_6; // @[CGRA.scala 200:20]
  wire [31:0] pes_15_io_in_7; // @[CGRA.scala 200:20]
  wire [31:0] pes_15_io_out_0; // @[CGRA.scala 200:20]
  wire  pes_16_clock; // @[CGRA.scala 200:20]
  wire  pes_16_reset; // @[CGRA.scala 200:20]
  wire  pes_16_io_cfg_en; // @[CGRA.scala 200:20]
  wire [11:0] pes_16_io_cfg_addr; // @[CGRA.scala 200:20]
  wire [31:0] pes_16_io_cfg_data; // @[CGRA.scala 200:20]
  wire  pes_16_io_en; // @[CGRA.scala 200:20]
  wire [31:0] pes_16_io_in_0; // @[CGRA.scala 200:20]
  wire [31:0] pes_16_io_in_1; // @[CGRA.scala 200:20]
  wire [31:0] pes_16_io_in_2; // @[CGRA.scala 200:20]
  wire [31:0] pes_16_io_in_3; // @[CGRA.scala 200:20]
  wire [31:0] pes_16_io_in_4; // @[CGRA.scala 200:20]
  wire [31:0] pes_16_io_in_5; // @[CGRA.scala 200:20]
  wire [31:0] pes_16_io_in_6; // @[CGRA.scala 200:20]
  wire [31:0] pes_16_io_in_7; // @[CGRA.scala 200:20]
  wire [31:0] pes_16_io_out_0; // @[CGRA.scala 200:20]
  wire  pes_17_clock; // @[CGRA.scala 200:20]
  wire  pes_17_reset; // @[CGRA.scala 200:20]
  wire  pes_17_io_cfg_en; // @[CGRA.scala 200:20]
  wire [11:0] pes_17_io_cfg_addr; // @[CGRA.scala 200:20]
  wire [31:0] pes_17_io_cfg_data; // @[CGRA.scala 200:20]
  wire  pes_17_io_en; // @[CGRA.scala 200:20]
  wire [31:0] pes_17_io_in_0; // @[CGRA.scala 200:20]
  wire [31:0] pes_17_io_in_1; // @[CGRA.scala 200:20]
  wire [31:0] pes_17_io_in_2; // @[CGRA.scala 200:20]
  wire [31:0] pes_17_io_in_3; // @[CGRA.scala 200:20]
  wire [31:0] pes_17_io_in_4; // @[CGRA.scala 200:20]
  wire [31:0] pes_17_io_in_5; // @[CGRA.scala 200:20]
  wire [31:0] pes_17_io_in_6; // @[CGRA.scala 200:20]
  wire [31:0] pes_17_io_in_7; // @[CGRA.scala 200:20]
  wire [31:0] pes_17_io_out_0; // @[CGRA.scala 200:20]
  wire  pes_18_clock; // @[CGRA.scala 200:20]
  wire  pes_18_reset; // @[CGRA.scala 200:20]
  wire  pes_18_io_cfg_en; // @[CGRA.scala 200:20]
  wire [11:0] pes_18_io_cfg_addr; // @[CGRA.scala 200:20]
  wire [31:0] pes_18_io_cfg_data; // @[CGRA.scala 200:20]
  wire  pes_18_io_en; // @[CGRA.scala 200:20]
  wire [31:0] pes_18_io_in_0; // @[CGRA.scala 200:20]
  wire [31:0] pes_18_io_in_1; // @[CGRA.scala 200:20]
  wire [31:0] pes_18_io_in_2; // @[CGRA.scala 200:20]
  wire [31:0] pes_18_io_in_3; // @[CGRA.scala 200:20]
  wire [31:0] pes_18_io_in_4; // @[CGRA.scala 200:20]
  wire [31:0] pes_18_io_in_5; // @[CGRA.scala 200:20]
  wire [31:0] pes_18_io_in_6; // @[CGRA.scala 200:20]
  wire [31:0] pes_18_io_in_7; // @[CGRA.scala 200:20]
  wire [31:0] pes_18_io_out_0; // @[CGRA.scala 200:20]
  wire  pes_19_clock; // @[CGRA.scala 200:20]
  wire  pes_19_reset; // @[CGRA.scala 200:20]
  wire  pes_19_io_cfg_en; // @[CGRA.scala 200:20]
  wire [11:0] pes_19_io_cfg_addr; // @[CGRA.scala 200:20]
  wire [31:0] pes_19_io_cfg_data; // @[CGRA.scala 200:20]
  wire  pes_19_io_en; // @[CGRA.scala 200:20]
  wire [31:0] pes_19_io_in_0; // @[CGRA.scala 200:20]
  wire [31:0] pes_19_io_in_1; // @[CGRA.scala 200:20]
  wire [31:0] pes_19_io_in_2; // @[CGRA.scala 200:20]
  wire [31:0] pes_19_io_in_3; // @[CGRA.scala 200:20]
  wire [31:0] pes_19_io_in_4; // @[CGRA.scala 200:20]
  wire [31:0] pes_19_io_in_5; // @[CGRA.scala 200:20]
  wire [31:0] pes_19_io_in_6; // @[CGRA.scala 200:20]
  wire [31:0] pes_19_io_in_7; // @[CGRA.scala 200:20]
  wire [31:0] pes_19_io_out_0; // @[CGRA.scala 200:20]
  wire  pes_20_clock; // @[CGRA.scala 200:20]
  wire  pes_20_reset; // @[CGRA.scala 200:20]
  wire  pes_20_io_cfg_en; // @[CGRA.scala 200:20]
  wire [11:0] pes_20_io_cfg_addr; // @[CGRA.scala 200:20]
  wire [31:0] pes_20_io_cfg_data; // @[CGRA.scala 200:20]
  wire  pes_20_io_en; // @[CGRA.scala 200:20]
  wire [31:0] pes_20_io_in_0; // @[CGRA.scala 200:20]
  wire [31:0] pes_20_io_in_1; // @[CGRA.scala 200:20]
  wire [31:0] pes_20_io_in_2; // @[CGRA.scala 200:20]
  wire [31:0] pes_20_io_in_3; // @[CGRA.scala 200:20]
  wire [31:0] pes_20_io_in_4; // @[CGRA.scala 200:20]
  wire [31:0] pes_20_io_in_5; // @[CGRA.scala 200:20]
  wire [31:0] pes_20_io_in_6; // @[CGRA.scala 200:20]
  wire [31:0] pes_20_io_in_7; // @[CGRA.scala 200:20]
  wire [31:0] pes_20_io_out_0; // @[CGRA.scala 200:20]
  wire  pes_21_clock; // @[CGRA.scala 200:20]
  wire  pes_21_reset; // @[CGRA.scala 200:20]
  wire  pes_21_io_cfg_en; // @[CGRA.scala 200:20]
  wire [11:0] pes_21_io_cfg_addr; // @[CGRA.scala 200:20]
  wire [31:0] pes_21_io_cfg_data; // @[CGRA.scala 200:20]
  wire  pes_21_io_en; // @[CGRA.scala 200:20]
  wire [31:0] pes_21_io_in_0; // @[CGRA.scala 200:20]
  wire [31:0] pes_21_io_in_1; // @[CGRA.scala 200:20]
  wire [31:0] pes_21_io_in_2; // @[CGRA.scala 200:20]
  wire [31:0] pes_21_io_in_3; // @[CGRA.scala 200:20]
  wire [31:0] pes_21_io_in_4; // @[CGRA.scala 200:20]
  wire [31:0] pes_21_io_in_5; // @[CGRA.scala 200:20]
  wire [31:0] pes_21_io_in_6; // @[CGRA.scala 200:20]
  wire [31:0] pes_21_io_in_7; // @[CGRA.scala 200:20]
  wire [31:0] pes_21_io_out_0; // @[CGRA.scala 200:20]
  wire  pes_22_clock; // @[CGRA.scala 200:20]
  wire  pes_22_reset; // @[CGRA.scala 200:20]
  wire  pes_22_io_cfg_en; // @[CGRA.scala 200:20]
  wire [11:0] pes_22_io_cfg_addr; // @[CGRA.scala 200:20]
  wire [31:0] pes_22_io_cfg_data; // @[CGRA.scala 200:20]
  wire  pes_22_io_en; // @[CGRA.scala 200:20]
  wire [31:0] pes_22_io_in_0; // @[CGRA.scala 200:20]
  wire [31:0] pes_22_io_in_1; // @[CGRA.scala 200:20]
  wire [31:0] pes_22_io_in_2; // @[CGRA.scala 200:20]
  wire [31:0] pes_22_io_in_3; // @[CGRA.scala 200:20]
  wire [31:0] pes_22_io_in_4; // @[CGRA.scala 200:20]
  wire [31:0] pes_22_io_in_5; // @[CGRA.scala 200:20]
  wire [31:0] pes_22_io_in_6; // @[CGRA.scala 200:20]
  wire [31:0] pes_22_io_in_7; // @[CGRA.scala 200:20]
  wire [31:0] pes_22_io_out_0; // @[CGRA.scala 200:20]
  wire  pes_23_clock; // @[CGRA.scala 200:20]
  wire  pes_23_reset; // @[CGRA.scala 200:20]
  wire  pes_23_io_cfg_en; // @[CGRA.scala 200:20]
  wire [11:0] pes_23_io_cfg_addr; // @[CGRA.scala 200:20]
  wire [31:0] pes_23_io_cfg_data; // @[CGRA.scala 200:20]
  wire  pes_23_io_en; // @[CGRA.scala 200:20]
  wire [31:0] pes_23_io_in_0; // @[CGRA.scala 200:20]
  wire [31:0] pes_23_io_in_1; // @[CGRA.scala 200:20]
  wire [31:0] pes_23_io_in_2; // @[CGRA.scala 200:20]
  wire [31:0] pes_23_io_in_3; // @[CGRA.scala 200:20]
  wire [31:0] pes_23_io_in_4; // @[CGRA.scala 200:20]
  wire [31:0] pes_23_io_in_5; // @[CGRA.scala 200:20]
  wire [31:0] pes_23_io_in_6; // @[CGRA.scala 200:20]
  wire [31:0] pes_23_io_in_7; // @[CGRA.scala 200:20]
  wire [31:0] pes_23_io_out_0; // @[CGRA.scala 200:20]
  wire  pes_24_clock; // @[CGRA.scala 200:20]
  wire  pes_24_reset; // @[CGRA.scala 200:20]
  wire  pes_24_io_cfg_en; // @[CGRA.scala 200:20]
  wire [11:0] pes_24_io_cfg_addr; // @[CGRA.scala 200:20]
  wire [31:0] pes_24_io_cfg_data; // @[CGRA.scala 200:20]
  wire  pes_24_io_en; // @[CGRA.scala 200:20]
  wire [31:0] pes_24_io_in_0; // @[CGRA.scala 200:20]
  wire [31:0] pes_24_io_in_1; // @[CGRA.scala 200:20]
  wire [31:0] pes_24_io_in_2; // @[CGRA.scala 200:20]
  wire [31:0] pes_24_io_in_3; // @[CGRA.scala 200:20]
  wire [31:0] pes_24_io_in_4; // @[CGRA.scala 200:20]
  wire [31:0] pes_24_io_in_5; // @[CGRA.scala 200:20]
  wire [31:0] pes_24_io_in_6; // @[CGRA.scala 200:20]
  wire [31:0] pes_24_io_in_7; // @[CGRA.scala 200:20]
  wire [31:0] pes_24_io_out_0; // @[CGRA.scala 200:20]
  wire  pes_25_clock; // @[CGRA.scala 200:20]
  wire  pes_25_reset; // @[CGRA.scala 200:20]
  wire  pes_25_io_cfg_en; // @[CGRA.scala 200:20]
  wire [11:0] pes_25_io_cfg_addr; // @[CGRA.scala 200:20]
  wire [31:0] pes_25_io_cfg_data; // @[CGRA.scala 200:20]
  wire  pes_25_io_en; // @[CGRA.scala 200:20]
  wire [31:0] pes_25_io_in_0; // @[CGRA.scala 200:20]
  wire [31:0] pes_25_io_in_1; // @[CGRA.scala 200:20]
  wire [31:0] pes_25_io_in_2; // @[CGRA.scala 200:20]
  wire [31:0] pes_25_io_in_3; // @[CGRA.scala 200:20]
  wire [31:0] pes_25_io_in_4; // @[CGRA.scala 200:20]
  wire [31:0] pes_25_io_in_5; // @[CGRA.scala 200:20]
  wire [31:0] pes_25_io_in_6; // @[CGRA.scala 200:20]
  wire [31:0] pes_25_io_in_7; // @[CGRA.scala 200:20]
  wire [31:0] pes_25_io_out_0; // @[CGRA.scala 200:20]
  wire  pes_26_clock; // @[CGRA.scala 200:20]
  wire  pes_26_reset; // @[CGRA.scala 200:20]
  wire  pes_26_io_cfg_en; // @[CGRA.scala 200:20]
  wire [11:0] pes_26_io_cfg_addr; // @[CGRA.scala 200:20]
  wire [31:0] pes_26_io_cfg_data; // @[CGRA.scala 200:20]
  wire  pes_26_io_en; // @[CGRA.scala 200:20]
  wire [31:0] pes_26_io_in_0; // @[CGRA.scala 200:20]
  wire [31:0] pes_26_io_in_1; // @[CGRA.scala 200:20]
  wire [31:0] pes_26_io_in_2; // @[CGRA.scala 200:20]
  wire [31:0] pes_26_io_in_3; // @[CGRA.scala 200:20]
  wire [31:0] pes_26_io_in_4; // @[CGRA.scala 200:20]
  wire [31:0] pes_26_io_in_5; // @[CGRA.scala 200:20]
  wire [31:0] pes_26_io_in_6; // @[CGRA.scala 200:20]
  wire [31:0] pes_26_io_in_7; // @[CGRA.scala 200:20]
  wire [31:0] pes_26_io_out_0; // @[CGRA.scala 200:20]
  wire  pes_27_clock; // @[CGRA.scala 200:20]
  wire  pes_27_reset; // @[CGRA.scala 200:20]
  wire  pes_27_io_cfg_en; // @[CGRA.scala 200:20]
  wire [11:0] pes_27_io_cfg_addr; // @[CGRA.scala 200:20]
  wire [31:0] pes_27_io_cfg_data; // @[CGRA.scala 200:20]
  wire  pes_27_io_en; // @[CGRA.scala 200:20]
  wire [31:0] pes_27_io_in_0; // @[CGRA.scala 200:20]
  wire [31:0] pes_27_io_in_1; // @[CGRA.scala 200:20]
  wire [31:0] pes_27_io_in_2; // @[CGRA.scala 200:20]
  wire [31:0] pes_27_io_in_3; // @[CGRA.scala 200:20]
  wire [31:0] pes_27_io_in_4; // @[CGRA.scala 200:20]
  wire [31:0] pes_27_io_in_5; // @[CGRA.scala 200:20]
  wire [31:0] pes_27_io_in_6; // @[CGRA.scala 200:20]
  wire [31:0] pes_27_io_in_7; // @[CGRA.scala 200:20]
  wire [31:0] pes_27_io_out_0; // @[CGRA.scala 200:20]
  wire  pes_28_clock; // @[CGRA.scala 200:20]
  wire  pes_28_reset; // @[CGRA.scala 200:20]
  wire  pes_28_io_cfg_en; // @[CGRA.scala 200:20]
  wire [11:0] pes_28_io_cfg_addr; // @[CGRA.scala 200:20]
  wire [31:0] pes_28_io_cfg_data; // @[CGRA.scala 200:20]
  wire  pes_28_io_en; // @[CGRA.scala 200:20]
  wire [31:0] pes_28_io_in_0; // @[CGRA.scala 200:20]
  wire [31:0] pes_28_io_in_1; // @[CGRA.scala 200:20]
  wire [31:0] pes_28_io_in_2; // @[CGRA.scala 200:20]
  wire [31:0] pes_28_io_in_3; // @[CGRA.scala 200:20]
  wire [31:0] pes_28_io_in_4; // @[CGRA.scala 200:20]
  wire [31:0] pes_28_io_in_5; // @[CGRA.scala 200:20]
  wire [31:0] pes_28_io_in_6; // @[CGRA.scala 200:20]
  wire [31:0] pes_28_io_in_7; // @[CGRA.scala 200:20]
  wire [31:0] pes_28_io_out_0; // @[CGRA.scala 200:20]
  wire  pes_29_clock; // @[CGRA.scala 200:20]
  wire  pes_29_reset; // @[CGRA.scala 200:20]
  wire  pes_29_io_cfg_en; // @[CGRA.scala 200:20]
  wire [11:0] pes_29_io_cfg_addr; // @[CGRA.scala 200:20]
  wire [31:0] pes_29_io_cfg_data; // @[CGRA.scala 200:20]
  wire  pes_29_io_en; // @[CGRA.scala 200:20]
  wire [31:0] pes_29_io_in_0; // @[CGRA.scala 200:20]
  wire [31:0] pes_29_io_in_1; // @[CGRA.scala 200:20]
  wire [31:0] pes_29_io_in_2; // @[CGRA.scala 200:20]
  wire [31:0] pes_29_io_in_3; // @[CGRA.scala 200:20]
  wire [31:0] pes_29_io_in_4; // @[CGRA.scala 200:20]
  wire [31:0] pes_29_io_in_5; // @[CGRA.scala 200:20]
  wire [31:0] pes_29_io_in_6; // @[CGRA.scala 200:20]
  wire [31:0] pes_29_io_in_7; // @[CGRA.scala 200:20]
  wire [31:0] pes_29_io_out_0; // @[CGRA.scala 200:20]
  wire  pes_30_clock; // @[CGRA.scala 200:20]
  wire  pes_30_reset; // @[CGRA.scala 200:20]
  wire  pes_30_io_cfg_en; // @[CGRA.scala 200:20]
  wire [11:0] pes_30_io_cfg_addr; // @[CGRA.scala 200:20]
  wire [31:0] pes_30_io_cfg_data; // @[CGRA.scala 200:20]
  wire  pes_30_io_en; // @[CGRA.scala 200:20]
  wire [31:0] pes_30_io_in_0; // @[CGRA.scala 200:20]
  wire [31:0] pes_30_io_in_1; // @[CGRA.scala 200:20]
  wire [31:0] pes_30_io_in_2; // @[CGRA.scala 200:20]
  wire [31:0] pes_30_io_in_3; // @[CGRA.scala 200:20]
  wire [31:0] pes_30_io_in_4; // @[CGRA.scala 200:20]
  wire [31:0] pes_30_io_in_5; // @[CGRA.scala 200:20]
  wire [31:0] pes_30_io_in_6; // @[CGRA.scala 200:20]
  wire [31:0] pes_30_io_in_7; // @[CGRA.scala 200:20]
  wire [31:0] pes_30_io_out_0; // @[CGRA.scala 200:20]
  wire  pes_31_clock; // @[CGRA.scala 200:20]
  wire  pes_31_reset; // @[CGRA.scala 200:20]
  wire  pes_31_io_cfg_en; // @[CGRA.scala 200:20]
  wire [11:0] pes_31_io_cfg_addr; // @[CGRA.scala 200:20]
  wire [31:0] pes_31_io_cfg_data; // @[CGRA.scala 200:20]
  wire  pes_31_io_en; // @[CGRA.scala 200:20]
  wire [31:0] pes_31_io_in_0; // @[CGRA.scala 200:20]
  wire [31:0] pes_31_io_in_1; // @[CGRA.scala 200:20]
  wire [31:0] pes_31_io_in_2; // @[CGRA.scala 200:20]
  wire [31:0] pes_31_io_in_3; // @[CGRA.scala 200:20]
  wire [31:0] pes_31_io_in_4; // @[CGRA.scala 200:20]
  wire [31:0] pes_31_io_in_5; // @[CGRA.scala 200:20]
  wire [31:0] pes_31_io_in_6; // @[CGRA.scala 200:20]
  wire [31:0] pes_31_io_in_7; // @[CGRA.scala 200:20]
  wire [31:0] pes_31_io_out_0; // @[CGRA.scala 200:20]
  wire  pes_32_clock; // @[CGRA.scala 200:20]
  wire  pes_32_reset; // @[CGRA.scala 200:20]
  wire  pes_32_io_cfg_en; // @[CGRA.scala 200:20]
  wire [11:0] pes_32_io_cfg_addr; // @[CGRA.scala 200:20]
  wire [31:0] pes_32_io_cfg_data; // @[CGRA.scala 200:20]
  wire  pes_32_io_en; // @[CGRA.scala 200:20]
  wire [31:0] pes_32_io_in_0; // @[CGRA.scala 200:20]
  wire [31:0] pes_32_io_in_1; // @[CGRA.scala 200:20]
  wire [31:0] pes_32_io_in_2; // @[CGRA.scala 200:20]
  wire [31:0] pes_32_io_in_3; // @[CGRA.scala 200:20]
  wire [31:0] pes_32_io_in_4; // @[CGRA.scala 200:20]
  wire [31:0] pes_32_io_in_5; // @[CGRA.scala 200:20]
  wire [31:0] pes_32_io_in_6; // @[CGRA.scala 200:20]
  wire [31:0] pes_32_io_in_7; // @[CGRA.scala 200:20]
  wire [31:0] pes_32_io_out_0; // @[CGRA.scala 200:20]
  wire  pes_33_clock; // @[CGRA.scala 200:20]
  wire  pes_33_reset; // @[CGRA.scala 200:20]
  wire  pes_33_io_cfg_en; // @[CGRA.scala 200:20]
  wire [11:0] pes_33_io_cfg_addr; // @[CGRA.scala 200:20]
  wire [31:0] pes_33_io_cfg_data; // @[CGRA.scala 200:20]
  wire  pes_33_io_en; // @[CGRA.scala 200:20]
  wire [31:0] pes_33_io_in_0; // @[CGRA.scala 200:20]
  wire [31:0] pes_33_io_in_1; // @[CGRA.scala 200:20]
  wire [31:0] pes_33_io_in_2; // @[CGRA.scala 200:20]
  wire [31:0] pes_33_io_in_3; // @[CGRA.scala 200:20]
  wire [31:0] pes_33_io_in_4; // @[CGRA.scala 200:20]
  wire [31:0] pes_33_io_in_5; // @[CGRA.scala 200:20]
  wire [31:0] pes_33_io_in_6; // @[CGRA.scala 200:20]
  wire [31:0] pes_33_io_in_7; // @[CGRA.scala 200:20]
  wire [31:0] pes_33_io_out_0; // @[CGRA.scala 200:20]
  wire  pes_34_clock; // @[CGRA.scala 200:20]
  wire  pes_34_reset; // @[CGRA.scala 200:20]
  wire  pes_34_io_cfg_en; // @[CGRA.scala 200:20]
  wire [11:0] pes_34_io_cfg_addr; // @[CGRA.scala 200:20]
  wire [31:0] pes_34_io_cfg_data; // @[CGRA.scala 200:20]
  wire  pes_34_io_en; // @[CGRA.scala 200:20]
  wire [31:0] pes_34_io_in_0; // @[CGRA.scala 200:20]
  wire [31:0] pes_34_io_in_1; // @[CGRA.scala 200:20]
  wire [31:0] pes_34_io_in_2; // @[CGRA.scala 200:20]
  wire [31:0] pes_34_io_in_3; // @[CGRA.scala 200:20]
  wire [31:0] pes_34_io_in_4; // @[CGRA.scala 200:20]
  wire [31:0] pes_34_io_in_5; // @[CGRA.scala 200:20]
  wire [31:0] pes_34_io_in_6; // @[CGRA.scala 200:20]
  wire [31:0] pes_34_io_in_7; // @[CGRA.scala 200:20]
  wire [31:0] pes_34_io_out_0; // @[CGRA.scala 200:20]
  wire  pes_35_clock; // @[CGRA.scala 200:20]
  wire  pes_35_reset; // @[CGRA.scala 200:20]
  wire  pes_35_io_cfg_en; // @[CGRA.scala 200:20]
  wire [11:0] pes_35_io_cfg_addr; // @[CGRA.scala 200:20]
  wire [31:0] pes_35_io_cfg_data; // @[CGRA.scala 200:20]
  wire  pes_35_io_en; // @[CGRA.scala 200:20]
  wire [31:0] pes_35_io_in_0; // @[CGRA.scala 200:20]
  wire [31:0] pes_35_io_in_1; // @[CGRA.scala 200:20]
  wire [31:0] pes_35_io_in_2; // @[CGRA.scala 200:20]
  wire [31:0] pes_35_io_in_3; // @[CGRA.scala 200:20]
  wire [31:0] pes_35_io_in_4; // @[CGRA.scala 200:20]
  wire [31:0] pes_35_io_in_5; // @[CGRA.scala 200:20]
  wire [31:0] pes_35_io_in_6; // @[CGRA.scala 200:20]
  wire [31:0] pes_35_io_in_7; // @[CGRA.scala 200:20]
  wire [31:0] pes_35_io_out_0; // @[CGRA.scala 200:20]
  wire  pes_36_clock; // @[CGRA.scala 200:20]
  wire  pes_36_reset; // @[CGRA.scala 200:20]
  wire  pes_36_io_cfg_en; // @[CGRA.scala 200:20]
  wire [11:0] pes_36_io_cfg_addr; // @[CGRA.scala 200:20]
  wire [31:0] pes_36_io_cfg_data; // @[CGRA.scala 200:20]
  wire  pes_36_io_en; // @[CGRA.scala 200:20]
  wire [31:0] pes_36_io_in_0; // @[CGRA.scala 200:20]
  wire [31:0] pes_36_io_in_1; // @[CGRA.scala 200:20]
  wire [31:0] pes_36_io_in_2; // @[CGRA.scala 200:20]
  wire [31:0] pes_36_io_in_3; // @[CGRA.scala 200:20]
  wire [31:0] pes_36_io_in_4; // @[CGRA.scala 200:20]
  wire [31:0] pes_36_io_in_5; // @[CGRA.scala 200:20]
  wire [31:0] pes_36_io_in_6; // @[CGRA.scala 200:20]
  wire [31:0] pes_36_io_in_7; // @[CGRA.scala 200:20]
  wire [31:0] pes_36_io_out_0; // @[CGRA.scala 200:20]
  wire  pes_37_clock; // @[CGRA.scala 200:20]
  wire  pes_37_reset; // @[CGRA.scala 200:20]
  wire  pes_37_io_cfg_en; // @[CGRA.scala 200:20]
  wire [11:0] pes_37_io_cfg_addr; // @[CGRA.scala 200:20]
  wire [31:0] pes_37_io_cfg_data; // @[CGRA.scala 200:20]
  wire  pes_37_io_en; // @[CGRA.scala 200:20]
  wire [31:0] pes_37_io_in_0; // @[CGRA.scala 200:20]
  wire [31:0] pes_37_io_in_1; // @[CGRA.scala 200:20]
  wire [31:0] pes_37_io_in_2; // @[CGRA.scala 200:20]
  wire [31:0] pes_37_io_in_3; // @[CGRA.scala 200:20]
  wire [31:0] pes_37_io_in_4; // @[CGRA.scala 200:20]
  wire [31:0] pes_37_io_in_5; // @[CGRA.scala 200:20]
  wire [31:0] pes_37_io_in_6; // @[CGRA.scala 200:20]
  wire [31:0] pes_37_io_in_7; // @[CGRA.scala 200:20]
  wire [31:0] pes_37_io_out_0; // @[CGRA.scala 200:20]
  wire  pes_38_clock; // @[CGRA.scala 200:20]
  wire  pes_38_reset; // @[CGRA.scala 200:20]
  wire  pes_38_io_cfg_en; // @[CGRA.scala 200:20]
  wire [11:0] pes_38_io_cfg_addr; // @[CGRA.scala 200:20]
  wire [31:0] pes_38_io_cfg_data; // @[CGRA.scala 200:20]
  wire  pes_38_io_en; // @[CGRA.scala 200:20]
  wire [31:0] pes_38_io_in_0; // @[CGRA.scala 200:20]
  wire [31:0] pes_38_io_in_1; // @[CGRA.scala 200:20]
  wire [31:0] pes_38_io_in_2; // @[CGRA.scala 200:20]
  wire [31:0] pes_38_io_in_3; // @[CGRA.scala 200:20]
  wire [31:0] pes_38_io_in_4; // @[CGRA.scala 200:20]
  wire [31:0] pes_38_io_in_5; // @[CGRA.scala 200:20]
  wire [31:0] pes_38_io_in_6; // @[CGRA.scala 200:20]
  wire [31:0] pes_38_io_in_7; // @[CGRA.scala 200:20]
  wire [31:0] pes_38_io_out_0; // @[CGRA.scala 200:20]
  wire  pes_39_clock; // @[CGRA.scala 200:20]
  wire  pes_39_reset; // @[CGRA.scala 200:20]
  wire  pes_39_io_cfg_en; // @[CGRA.scala 200:20]
  wire [11:0] pes_39_io_cfg_addr; // @[CGRA.scala 200:20]
  wire [31:0] pes_39_io_cfg_data; // @[CGRA.scala 200:20]
  wire  pes_39_io_en; // @[CGRA.scala 200:20]
  wire [31:0] pes_39_io_in_0; // @[CGRA.scala 200:20]
  wire [31:0] pes_39_io_in_1; // @[CGRA.scala 200:20]
  wire [31:0] pes_39_io_in_2; // @[CGRA.scala 200:20]
  wire [31:0] pes_39_io_in_3; // @[CGRA.scala 200:20]
  wire [31:0] pes_39_io_in_4; // @[CGRA.scala 200:20]
  wire [31:0] pes_39_io_in_5; // @[CGRA.scala 200:20]
  wire [31:0] pes_39_io_in_6; // @[CGRA.scala 200:20]
  wire [31:0] pes_39_io_in_7; // @[CGRA.scala 200:20]
  wire [31:0] pes_39_io_out_0; // @[CGRA.scala 200:20]
  wire  pes_40_clock; // @[CGRA.scala 200:20]
  wire  pes_40_reset; // @[CGRA.scala 200:20]
  wire  pes_40_io_cfg_en; // @[CGRA.scala 200:20]
  wire [11:0] pes_40_io_cfg_addr; // @[CGRA.scala 200:20]
  wire [31:0] pes_40_io_cfg_data; // @[CGRA.scala 200:20]
  wire  pes_40_io_en; // @[CGRA.scala 200:20]
  wire [31:0] pes_40_io_in_0; // @[CGRA.scala 200:20]
  wire [31:0] pes_40_io_in_1; // @[CGRA.scala 200:20]
  wire [31:0] pes_40_io_in_2; // @[CGRA.scala 200:20]
  wire [31:0] pes_40_io_in_3; // @[CGRA.scala 200:20]
  wire [31:0] pes_40_io_in_4; // @[CGRA.scala 200:20]
  wire [31:0] pes_40_io_in_5; // @[CGRA.scala 200:20]
  wire [31:0] pes_40_io_in_6; // @[CGRA.scala 200:20]
  wire [31:0] pes_40_io_in_7; // @[CGRA.scala 200:20]
  wire [31:0] pes_40_io_out_0; // @[CGRA.scala 200:20]
  wire  pes_41_clock; // @[CGRA.scala 200:20]
  wire  pes_41_reset; // @[CGRA.scala 200:20]
  wire  pes_41_io_cfg_en; // @[CGRA.scala 200:20]
  wire [11:0] pes_41_io_cfg_addr; // @[CGRA.scala 200:20]
  wire [31:0] pes_41_io_cfg_data; // @[CGRA.scala 200:20]
  wire  pes_41_io_en; // @[CGRA.scala 200:20]
  wire [31:0] pes_41_io_in_0; // @[CGRA.scala 200:20]
  wire [31:0] pes_41_io_in_1; // @[CGRA.scala 200:20]
  wire [31:0] pes_41_io_in_2; // @[CGRA.scala 200:20]
  wire [31:0] pes_41_io_in_3; // @[CGRA.scala 200:20]
  wire [31:0] pes_41_io_in_4; // @[CGRA.scala 200:20]
  wire [31:0] pes_41_io_in_5; // @[CGRA.scala 200:20]
  wire [31:0] pes_41_io_in_6; // @[CGRA.scala 200:20]
  wire [31:0] pes_41_io_in_7; // @[CGRA.scala 200:20]
  wire [31:0] pes_41_io_out_0; // @[CGRA.scala 200:20]
  wire  pes_42_clock; // @[CGRA.scala 200:20]
  wire  pes_42_reset; // @[CGRA.scala 200:20]
  wire  pes_42_io_cfg_en; // @[CGRA.scala 200:20]
  wire [11:0] pes_42_io_cfg_addr; // @[CGRA.scala 200:20]
  wire [31:0] pes_42_io_cfg_data; // @[CGRA.scala 200:20]
  wire  pes_42_io_en; // @[CGRA.scala 200:20]
  wire [31:0] pes_42_io_in_0; // @[CGRA.scala 200:20]
  wire [31:0] pes_42_io_in_1; // @[CGRA.scala 200:20]
  wire [31:0] pes_42_io_in_2; // @[CGRA.scala 200:20]
  wire [31:0] pes_42_io_in_3; // @[CGRA.scala 200:20]
  wire [31:0] pes_42_io_in_4; // @[CGRA.scala 200:20]
  wire [31:0] pes_42_io_in_5; // @[CGRA.scala 200:20]
  wire [31:0] pes_42_io_in_6; // @[CGRA.scala 200:20]
  wire [31:0] pes_42_io_in_7; // @[CGRA.scala 200:20]
  wire [31:0] pes_42_io_out_0; // @[CGRA.scala 200:20]
  wire  pes_43_clock; // @[CGRA.scala 200:20]
  wire  pes_43_reset; // @[CGRA.scala 200:20]
  wire  pes_43_io_cfg_en; // @[CGRA.scala 200:20]
  wire [11:0] pes_43_io_cfg_addr; // @[CGRA.scala 200:20]
  wire [31:0] pes_43_io_cfg_data; // @[CGRA.scala 200:20]
  wire  pes_43_io_en; // @[CGRA.scala 200:20]
  wire [31:0] pes_43_io_in_0; // @[CGRA.scala 200:20]
  wire [31:0] pes_43_io_in_1; // @[CGRA.scala 200:20]
  wire [31:0] pes_43_io_in_2; // @[CGRA.scala 200:20]
  wire [31:0] pes_43_io_in_3; // @[CGRA.scala 200:20]
  wire [31:0] pes_43_io_in_4; // @[CGRA.scala 200:20]
  wire [31:0] pes_43_io_in_5; // @[CGRA.scala 200:20]
  wire [31:0] pes_43_io_in_6; // @[CGRA.scala 200:20]
  wire [31:0] pes_43_io_in_7; // @[CGRA.scala 200:20]
  wire [31:0] pes_43_io_out_0; // @[CGRA.scala 200:20]
  wire  pes_44_clock; // @[CGRA.scala 200:20]
  wire  pes_44_reset; // @[CGRA.scala 200:20]
  wire  pes_44_io_cfg_en; // @[CGRA.scala 200:20]
  wire [11:0] pes_44_io_cfg_addr; // @[CGRA.scala 200:20]
  wire [31:0] pes_44_io_cfg_data; // @[CGRA.scala 200:20]
  wire  pes_44_io_en; // @[CGRA.scala 200:20]
  wire [31:0] pes_44_io_in_0; // @[CGRA.scala 200:20]
  wire [31:0] pes_44_io_in_1; // @[CGRA.scala 200:20]
  wire [31:0] pes_44_io_in_2; // @[CGRA.scala 200:20]
  wire [31:0] pes_44_io_in_3; // @[CGRA.scala 200:20]
  wire [31:0] pes_44_io_in_4; // @[CGRA.scala 200:20]
  wire [31:0] pes_44_io_in_5; // @[CGRA.scala 200:20]
  wire [31:0] pes_44_io_in_6; // @[CGRA.scala 200:20]
  wire [31:0] pes_44_io_in_7; // @[CGRA.scala 200:20]
  wire [31:0] pes_44_io_out_0; // @[CGRA.scala 200:20]
  wire  pes_45_clock; // @[CGRA.scala 200:20]
  wire  pes_45_reset; // @[CGRA.scala 200:20]
  wire  pes_45_io_cfg_en; // @[CGRA.scala 200:20]
  wire [11:0] pes_45_io_cfg_addr; // @[CGRA.scala 200:20]
  wire [31:0] pes_45_io_cfg_data; // @[CGRA.scala 200:20]
  wire  pes_45_io_en; // @[CGRA.scala 200:20]
  wire [31:0] pes_45_io_in_0; // @[CGRA.scala 200:20]
  wire [31:0] pes_45_io_in_1; // @[CGRA.scala 200:20]
  wire [31:0] pes_45_io_in_2; // @[CGRA.scala 200:20]
  wire [31:0] pes_45_io_in_3; // @[CGRA.scala 200:20]
  wire [31:0] pes_45_io_in_4; // @[CGRA.scala 200:20]
  wire [31:0] pes_45_io_in_5; // @[CGRA.scala 200:20]
  wire [31:0] pes_45_io_in_6; // @[CGRA.scala 200:20]
  wire [31:0] pes_45_io_in_7; // @[CGRA.scala 200:20]
  wire [31:0] pes_45_io_out_0; // @[CGRA.scala 200:20]
  wire  pes_46_clock; // @[CGRA.scala 200:20]
  wire  pes_46_reset; // @[CGRA.scala 200:20]
  wire  pes_46_io_cfg_en; // @[CGRA.scala 200:20]
  wire [11:0] pes_46_io_cfg_addr; // @[CGRA.scala 200:20]
  wire [31:0] pes_46_io_cfg_data; // @[CGRA.scala 200:20]
  wire  pes_46_io_en; // @[CGRA.scala 200:20]
  wire [31:0] pes_46_io_in_0; // @[CGRA.scala 200:20]
  wire [31:0] pes_46_io_in_1; // @[CGRA.scala 200:20]
  wire [31:0] pes_46_io_in_2; // @[CGRA.scala 200:20]
  wire [31:0] pes_46_io_in_3; // @[CGRA.scala 200:20]
  wire [31:0] pes_46_io_in_4; // @[CGRA.scala 200:20]
  wire [31:0] pes_46_io_in_5; // @[CGRA.scala 200:20]
  wire [31:0] pes_46_io_in_6; // @[CGRA.scala 200:20]
  wire [31:0] pes_46_io_in_7; // @[CGRA.scala 200:20]
  wire [31:0] pes_46_io_out_0; // @[CGRA.scala 200:20]
  wire  pes_47_clock; // @[CGRA.scala 200:20]
  wire  pes_47_reset; // @[CGRA.scala 200:20]
  wire  pes_47_io_cfg_en; // @[CGRA.scala 200:20]
  wire [11:0] pes_47_io_cfg_addr; // @[CGRA.scala 200:20]
  wire [31:0] pes_47_io_cfg_data; // @[CGRA.scala 200:20]
  wire  pes_47_io_en; // @[CGRA.scala 200:20]
  wire [31:0] pes_47_io_in_0; // @[CGRA.scala 200:20]
  wire [31:0] pes_47_io_in_1; // @[CGRA.scala 200:20]
  wire [31:0] pes_47_io_in_2; // @[CGRA.scala 200:20]
  wire [31:0] pes_47_io_in_3; // @[CGRA.scala 200:20]
  wire [31:0] pes_47_io_in_4; // @[CGRA.scala 200:20]
  wire [31:0] pes_47_io_in_5; // @[CGRA.scala 200:20]
  wire [31:0] pes_47_io_in_6; // @[CGRA.scala 200:20]
  wire [31:0] pes_47_io_in_7; // @[CGRA.scala 200:20]
  wire [31:0] pes_47_io_out_0; // @[CGRA.scala 200:20]
  wire  pes_48_clock; // @[CGRA.scala 200:20]
  wire  pes_48_reset; // @[CGRA.scala 200:20]
  wire  pes_48_io_cfg_en; // @[CGRA.scala 200:20]
  wire [11:0] pes_48_io_cfg_addr; // @[CGRA.scala 200:20]
  wire [31:0] pes_48_io_cfg_data; // @[CGRA.scala 200:20]
  wire  pes_48_io_en; // @[CGRA.scala 200:20]
  wire [31:0] pes_48_io_in_0; // @[CGRA.scala 200:20]
  wire [31:0] pes_48_io_in_1; // @[CGRA.scala 200:20]
  wire [31:0] pes_48_io_in_2; // @[CGRA.scala 200:20]
  wire [31:0] pes_48_io_in_3; // @[CGRA.scala 200:20]
  wire [31:0] pes_48_io_in_4; // @[CGRA.scala 200:20]
  wire [31:0] pes_48_io_in_5; // @[CGRA.scala 200:20]
  wire [31:0] pes_48_io_in_6; // @[CGRA.scala 200:20]
  wire [31:0] pes_48_io_in_7; // @[CGRA.scala 200:20]
  wire [31:0] pes_48_io_out_0; // @[CGRA.scala 200:20]
  wire  pes_49_clock; // @[CGRA.scala 200:20]
  wire  pes_49_reset; // @[CGRA.scala 200:20]
  wire  pes_49_io_cfg_en; // @[CGRA.scala 200:20]
  wire [11:0] pes_49_io_cfg_addr; // @[CGRA.scala 200:20]
  wire [31:0] pes_49_io_cfg_data; // @[CGRA.scala 200:20]
  wire  pes_49_io_en; // @[CGRA.scala 200:20]
  wire [31:0] pes_49_io_in_0; // @[CGRA.scala 200:20]
  wire [31:0] pes_49_io_in_1; // @[CGRA.scala 200:20]
  wire [31:0] pes_49_io_in_2; // @[CGRA.scala 200:20]
  wire [31:0] pes_49_io_in_3; // @[CGRA.scala 200:20]
  wire [31:0] pes_49_io_in_4; // @[CGRA.scala 200:20]
  wire [31:0] pes_49_io_in_5; // @[CGRA.scala 200:20]
  wire [31:0] pes_49_io_in_6; // @[CGRA.scala 200:20]
  wire [31:0] pes_49_io_in_7; // @[CGRA.scala 200:20]
  wire [31:0] pes_49_io_out_0; // @[CGRA.scala 200:20]
  wire  pes_50_clock; // @[CGRA.scala 200:20]
  wire  pes_50_reset; // @[CGRA.scala 200:20]
  wire  pes_50_io_cfg_en; // @[CGRA.scala 200:20]
  wire [11:0] pes_50_io_cfg_addr; // @[CGRA.scala 200:20]
  wire [31:0] pes_50_io_cfg_data; // @[CGRA.scala 200:20]
  wire  pes_50_io_en; // @[CGRA.scala 200:20]
  wire [31:0] pes_50_io_in_0; // @[CGRA.scala 200:20]
  wire [31:0] pes_50_io_in_1; // @[CGRA.scala 200:20]
  wire [31:0] pes_50_io_in_2; // @[CGRA.scala 200:20]
  wire [31:0] pes_50_io_in_3; // @[CGRA.scala 200:20]
  wire [31:0] pes_50_io_in_4; // @[CGRA.scala 200:20]
  wire [31:0] pes_50_io_in_5; // @[CGRA.scala 200:20]
  wire [31:0] pes_50_io_in_6; // @[CGRA.scala 200:20]
  wire [31:0] pes_50_io_in_7; // @[CGRA.scala 200:20]
  wire [31:0] pes_50_io_out_0; // @[CGRA.scala 200:20]
  wire  pes_51_clock; // @[CGRA.scala 200:20]
  wire  pes_51_reset; // @[CGRA.scala 200:20]
  wire  pes_51_io_cfg_en; // @[CGRA.scala 200:20]
  wire [11:0] pes_51_io_cfg_addr; // @[CGRA.scala 200:20]
  wire [31:0] pes_51_io_cfg_data; // @[CGRA.scala 200:20]
  wire  pes_51_io_en; // @[CGRA.scala 200:20]
  wire [31:0] pes_51_io_in_0; // @[CGRA.scala 200:20]
  wire [31:0] pes_51_io_in_1; // @[CGRA.scala 200:20]
  wire [31:0] pes_51_io_in_2; // @[CGRA.scala 200:20]
  wire [31:0] pes_51_io_in_3; // @[CGRA.scala 200:20]
  wire [31:0] pes_51_io_in_4; // @[CGRA.scala 200:20]
  wire [31:0] pes_51_io_in_5; // @[CGRA.scala 200:20]
  wire [31:0] pes_51_io_in_6; // @[CGRA.scala 200:20]
  wire [31:0] pes_51_io_in_7; // @[CGRA.scala 200:20]
  wire [31:0] pes_51_io_out_0; // @[CGRA.scala 200:20]
  wire  pes_52_clock; // @[CGRA.scala 200:20]
  wire  pes_52_reset; // @[CGRA.scala 200:20]
  wire  pes_52_io_cfg_en; // @[CGRA.scala 200:20]
  wire [11:0] pes_52_io_cfg_addr; // @[CGRA.scala 200:20]
  wire [31:0] pes_52_io_cfg_data; // @[CGRA.scala 200:20]
  wire  pes_52_io_en; // @[CGRA.scala 200:20]
  wire [31:0] pes_52_io_in_0; // @[CGRA.scala 200:20]
  wire [31:0] pes_52_io_in_1; // @[CGRA.scala 200:20]
  wire [31:0] pes_52_io_in_2; // @[CGRA.scala 200:20]
  wire [31:0] pes_52_io_in_3; // @[CGRA.scala 200:20]
  wire [31:0] pes_52_io_in_4; // @[CGRA.scala 200:20]
  wire [31:0] pes_52_io_in_5; // @[CGRA.scala 200:20]
  wire [31:0] pes_52_io_in_6; // @[CGRA.scala 200:20]
  wire [31:0] pes_52_io_in_7; // @[CGRA.scala 200:20]
  wire [31:0] pes_52_io_out_0; // @[CGRA.scala 200:20]
  wire  pes_53_clock; // @[CGRA.scala 200:20]
  wire  pes_53_reset; // @[CGRA.scala 200:20]
  wire  pes_53_io_cfg_en; // @[CGRA.scala 200:20]
  wire [11:0] pes_53_io_cfg_addr; // @[CGRA.scala 200:20]
  wire [31:0] pes_53_io_cfg_data; // @[CGRA.scala 200:20]
  wire  pes_53_io_en; // @[CGRA.scala 200:20]
  wire [31:0] pes_53_io_in_0; // @[CGRA.scala 200:20]
  wire [31:0] pes_53_io_in_1; // @[CGRA.scala 200:20]
  wire [31:0] pes_53_io_in_2; // @[CGRA.scala 200:20]
  wire [31:0] pes_53_io_in_3; // @[CGRA.scala 200:20]
  wire [31:0] pes_53_io_in_4; // @[CGRA.scala 200:20]
  wire [31:0] pes_53_io_in_5; // @[CGRA.scala 200:20]
  wire [31:0] pes_53_io_in_6; // @[CGRA.scala 200:20]
  wire [31:0] pes_53_io_in_7; // @[CGRA.scala 200:20]
  wire [31:0] pes_53_io_out_0; // @[CGRA.scala 200:20]
  wire  pes_54_clock; // @[CGRA.scala 200:20]
  wire  pes_54_reset; // @[CGRA.scala 200:20]
  wire  pes_54_io_cfg_en; // @[CGRA.scala 200:20]
  wire [11:0] pes_54_io_cfg_addr; // @[CGRA.scala 200:20]
  wire [31:0] pes_54_io_cfg_data; // @[CGRA.scala 200:20]
  wire  pes_54_io_en; // @[CGRA.scala 200:20]
  wire [31:0] pes_54_io_in_0; // @[CGRA.scala 200:20]
  wire [31:0] pes_54_io_in_1; // @[CGRA.scala 200:20]
  wire [31:0] pes_54_io_in_2; // @[CGRA.scala 200:20]
  wire [31:0] pes_54_io_in_3; // @[CGRA.scala 200:20]
  wire [31:0] pes_54_io_in_4; // @[CGRA.scala 200:20]
  wire [31:0] pes_54_io_in_5; // @[CGRA.scala 200:20]
  wire [31:0] pes_54_io_in_6; // @[CGRA.scala 200:20]
  wire [31:0] pes_54_io_in_7; // @[CGRA.scala 200:20]
  wire [31:0] pes_54_io_out_0; // @[CGRA.scala 200:20]
  wire  pes_55_clock; // @[CGRA.scala 200:20]
  wire  pes_55_reset; // @[CGRA.scala 200:20]
  wire  pes_55_io_cfg_en; // @[CGRA.scala 200:20]
  wire [11:0] pes_55_io_cfg_addr; // @[CGRA.scala 200:20]
  wire [31:0] pes_55_io_cfg_data; // @[CGRA.scala 200:20]
  wire  pes_55_io_en; // @[CGRA.scala 200:20]
  wire [31:0] pes_55_io_in_0; // @[CGRA.scala 200:20]
  wire [31:0] pes_55_io_in_1; // @[CGRA.scala 200:20]
  wire [31:0] pes_55_io_in_2; // @[CGRA.scala 200:20]
  wire [31:0] pes_55_io_in_3; // @[CGRA.scala 200:20]
  wire [31:0] pes_55_io_in_4; // @[CGRA.scala 200:20]
  wire [31:0] pes_55_io_in_5; // @[CGRA.scala 200:20]
  wire [31:0] pes_55_io_in_6; // @[CGRA.scala 200:20]
  wire [31:0] pes_55_io_in_7; // @[CGRA.scala 200:20]
  wire [31:0] pes_55_io_out_0; // @[CGRA.scala 200:20]
  wire  pes_56_clock; // @[CGRA.scala 200:20]
  wire  pes_56_reset; // @[CGRA.scala 200:20]
  wire  pes_56_io_cfg_en; // @[CGRA.scala 200:20]
  wire [11:0] pes_56_io_cfg_addr; // @[CGRA.scala 200:20]
  wire [31:0] pes_56_io_cfg_data; // @[CGRA.scala 200:20]
  wire  pes_56_io_en; // @[CGRA.scala 200:20]
  wire [31:0] pes_56_io_in_0; // @[CGRA.scala 200:20]
  wire [31:0] pes_56_io_in_1; // @[CGRA.scala 200:20]
  wire [31:0] pes_56_io_in_2; // @[CGRA.scala 200:20]
  wire [31:0] pes_56_io_in_3; // @[CGRA.scala 200:20]
  wire [31:0] pes_56_io_in_4; // @[CGRA.scala 200:20]
  wire [31:0] pes_56_io_in_5; // @[CGRA.scala 200:20]
  wire [31:0] pes_56_io_in_6; // @[CGRA.scala 200:20]
  wire [31:0] pes_56_io_in_7; // @[CGRA.scala 200:20]
  wire [31:0] pes_56_io_out_0; // @[CGRA.scala 200:20]
  wire  pes_57_clock; // @[CGRA.scala 200:20]
  wire  pes_57_reset; // @[CGRA.scala 200:20]
  wire  pes_57_io_cfg_en; // @[CGRA.scala 200:20]
  wire [11:0] pes_57_io_cfg_addr; // @[CGRA.scala 200:20]
  wire [31:0] pes_57_io_cfg_data; // @[CGRA.scala 200:20]
  wire  pes_57_io_en; // @[CGRA.scala 200:20]
  wire [31:0] pes_57_io_in_0; // @[CGRA.scala 200:20]
  wire [31:0] pes_57_io_in_1; // @[CGRA.scala 200:20]
  wire [31:0] pes_57_io_in_2; // @[CGRA.scala 200:20]
  wire [31:0] pes_57_io_in_3; // @[CGRA.scala 200:20]
  wire [31:0] pes_57_io_in_4; // @[CGRA.scala 200:20]
  wire [31:0] pes_57_io_in_5; // @[CGRA.scala 200:20]
  wire [31:0] pes_57_io_in_6; // @[CGRA.scala 200:20]
  wire [31:0] pes_57_io_in_7; // @[CGRA.scala 200:20]
  wire [31:0] pes_57_io_out_0; // @[CGRA.scala 200:20]
  wire  pes_58_clock; // @[CGRA.scala 200:20]
  wire  pes_58_reset; // @[CGRA.scala 200:20]
  wire  pes_58_io_cfg_en; // @[CGRA.scala 200:20]
  wire [11:0] pes_58_io_cfg_addr; // @[CGRA.scala 200:20]
  wire [31:0] pes_58_io_cfg_data; // @[CGRA.scala 200:20]
  wire  pes_58_io_en; // @[CGRA.scala 200:20]
  wire [31:0] pes_58_io_in_0; // @[CGRA.scala 200:20]
  wire [31:0] pes_58_io_in_1; // @[CGRA.scala 200:20]
  wire [31:0] pes_58_io_in_2; // @[CGRA.scala 200:20]
  wire [31:0] pes_58_io_in_3; // @[CGRA.scala 200:20]
  wire [31:0] pes_58_io_in_4; // @[CGRA.scala 200:20]
  wire [31:0] pes_58_io_in_5; // @[CGRA.scala 200:20]
  wire [31:0] pes_58_io_in_6; // @[CGRA.scala 200:20]
  wire [31:0] pes_58_io_in_7; // @[CGRA.scala 200:20]
  wire [31:0] pes_58_io_out_0; // @[CGRA.scala 200:20]
  wire  pes_59_clock; // @[CGRA.scala 200:20]
  wire  pes_59_reset; // @[CGRA.scala 200:20]
  wire  pes_59_io_cfg_en; // @[CGRA.scala 200:20]
  wire [11:0] pes_59_io_cfg_addr; // @[CGRA.scala 200:20]
  wire [31:0] pes_59_io_cfg_data; // @[CGRA.scala 200:20]
  wire  pes_59_io_en; // @[CGRA.scala 200:20]
  wire [31:0] pes_59_io_in_0; // @[CGRA.scala 200:20]
  wire [31:0] pes_59_io_in_1; // @[CGRA.scala 200:20]
  wire [31:0] pes_59_io_in_2; // @[CGRA.scala 200:20]
  wire [31:0] pes_59_io_in_3; // @[CGRA.scala 200:20]
  wire [31:0] pes_59_io_in_4; // @[CGRA.scala 200:20]
  wire [31:0] pes_59_io_in_5; // @[CGRA.scala 200:20]
  wire [31:0] pes_59_io_in_6; // @[CGRA.scala 200:20]
  wire [31:0] pes_59_io_in_7; // @[CGRA.scala 200:20]
  wire [31:0] pes_59_io_out_0; // @[CGRA.scala 200:20]
  wire  pes_60_clock; // @[CGRA.scala 200:20]
  wire  pes_60_reset; // @[CGRA.scala 200:20]
  wire  pes_60_io_cfg_en; // @[CGRA.scala 200:20]
  wire [11:0] pes_60_io_cfg_addr; // @[CGRA.scala 200:20]
  wire [31:0] pes_60_io_cfg_data; // @[CGRA.scala 200:20]
  wire  pes_60_io_en; // @[CGRA.scala 200:20]
  wire [31:0] pes_60_io_in_0; // @[CGRA.scala 200:20]
  wire [31:0] pes_60_io_in_1; // @[CGRA.scala 200:20]
  wire [31:0] pes_60_io_in_2; // @[CGRA.scala 200:20]
  wire [31:0] pes_60_io_in_3; // @[CGRA.scala 200:20]
  wire [31:0] pes_60_io_in_4; // @[CGRA.scala 200:20]
  wire [31:0] pes_60_io_in_5; // @[CGRA.scala 200:20]
  wire [31:0] pes_60_io_in_6; // @[CGRA.scala 200:20]
  wire [31:0] pes_60_io_in_7; // @[CGRA.scala 200:20]
  wire [31:0] pes_60_io_out_0; // @[CGRA.scala 200:20]
  wire  pes_61_clock; // @[CGRA.scala 200:20]
  wire  pes_61_reset; // @[CGRA.scala 200:20]
  wire  pes_61_io_cfg_en; // @[CGRA.scala 200:20]
  wire [11:0] pes_61_io_cfg_addr; // @[CGRA.scala 200:20]
  wire [31:0] pes_61_io_cfg_data; // @[CGRA.scala 200:20]
  wire  pes_61_io_en; // @[CGRA.scala 200:20]
  wire [31:0] pes_61_io_in_0; // @[CGRA.scala 200:20]
  wire [31:0] pes_61_io_in_1; // @[CGRA.scala 200:20]
  wire [31:0] pes_61_io_in_2; // @[CGRA.scala 200:20]
  wire [31:0] pes_61_io_in_3; // @[CGRA.scala 200:20]
  wire [31:0] pes_61_io_in_4; // @[CGRA.scala 200:20]
  wire [31:0] pes_61_io_in_5; // @[CGRA.scala 200:20]
  wire [31:0] pes_61_io_in_6; // @[CGRA.scala 200:20]
  wire [31:0] pes_61_io_in_7; // @[CGRA.scala 200:20]
  wire [31:0] pes_61_io_out_0; // @[CGRA.scala 200:20]
  wire  pes_62_clock; // @[CGRA.scala 200:20]
  wire  pes_62_reset; // @[CGRA.scala 200:20]
  wire  pes_62_io_cfg_en; // @[CGRA.scala 200:20]
  wire [11:0] pes_62_io_cfg_addr; // @[CGRA.scala 200:20]
  wire [31:0] pes_62_io_cfg_data; // @[CGRA.scala 200:20]
  wire  pes_62_io_en; // @[CGRA.scala 200:20]
  wire [31:0] pes_62_io_in_0; // @[CGRA.scala 200:20]
  wire [31:0] pes_62_io_in_1; // @[CGRA.scala 200:20]
  wire [31:0] pes_62_io_in_2; // @[CGRA.scala 200:20]
  wire [31:0] pes_62_io_in_3; // @[CGRA.scala 200:20]
  wire [31:0] pes_62_io_in_4; // @[CGRA.scala 200:20]
  wire [31:0] pes_62_io_in_5; // @[CGRA.scala 200:20]
  wire [31:0] pes_62_io_in_6; // @[CGRA.scala 200:20]
  wire [31:0] pes_62_io_in_7; // @[CGRA.scala 200:20]
  wire [31:0] pes_62_io_out_0; // @[CGRA.scala 200:20]
  wire  pes_63_clock; // @[CGRA.scala 200:20]
  wire  pes_63_reset; // @[CGRA.scala 200:20]
  wire  pes_63_io_cfg_en; // @[CGRA.scala 200:20]
  wire [11:0] pes_63_io_cfg_addr; // @[CGRA.scala 200:20]
  wire [31:0] pes_63_io_cfg_data; // @[CGRA.scala 200:20]
  wire  pes_63_io_en; // @[CGRA.scala 200:20]
  wire [31:0] pes_63_io_in_0; // @[CGRA.scala 200:20]
  wire [31:0] pes_63_io_in_1; // @[CGRA.scala 200:20]
  wire [31:0] pes_63_io_in_2; // @[CGRA.scala 200:20]
  wire [31:0] pes_63_io_in_3; // @[CGRA.scala 200:20]
  wire [31:0] pes_63_io_in_4; // @[CGRA.scala 200:20]
  wire [31:0] pes_63_io_in_5; // @[CGRA.scala 200:20]
  wire [31:0] pes_63_io_in_6; // @[CGRA.scala 200:20]
  wire [31:0] pes_63_io_in_7; // @[CGRA.scala 200:20]
  wire [31:0] pes_63_io_out_0; // @[CGRA.scala 200:20]
  wire  gibs_0_clock; // @[CGRA.scala 273:21]
  wire  gibs_0_reset; // @[CGRA.scala 273:21]
  wire  gibs_0_io_cfg_en; // @[CGRA.scala 273:21]
  wire [11:0] gibs_0_io_cfg_addr; // @[CGRA.scala 273:21]
  wire [31:0] gibs_0_io_cfg_data; // @[CGRA.scala 273:21]
  wire [31:0] gibs_0_io_ipinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_0_io_opinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_0_io_ipinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_0_io_ipinSE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_0_io_opinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_0_io_itrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_0_io_otrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_0_io_itrackS_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_0_io_otrackS_0; // @[CGRA.scala 273:21]
  wire  gibs_1_clock; // @[CGRA.scala 273:21]
  wire  gibs_1_reset; // @[CGRA.scala 273:21]
  wire  gibs_1_io_cfg_en; // @[CGRA.scala 273:21]
  wire [11:0] gibs_1_io_cfg_addr; // @[CGRA.scala 273:21]
  wire [31:0] gibs_1_io_cfg_data; // @[CGRA.scala 273:21]
  wire [31:0] gibs_1_io_ipinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_1_io_opinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_1_io_ipinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_1_io_opinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_1_io_ipinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_1_io_ipinSE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_1_io_opinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_1_io_ipinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_1_io_ipinSW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_1_io_opinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_1_io_itrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_1_io_otrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_1_io_itrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_1_io_otrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_1_io_itrackS_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_1_io_otrackS_0; // @[CGRA.scala 273:21]
  wire  gibs_2_clock; // @[CGRA.scala 273:21]
  wire  gibs_2_reset; // @[CGRA.scala 273:21]
  wire  gibs_2_io_cfg_en; // @[CGRA.scala 273:21]
  wire [11:0] gibs_2_io_cfg_addr; // @[CGRA.scala 273:21]
  wire [31:0] gibs_2_io_cfg_data; // @[CGRA.scala 273:21]
  wire [31:0] gibs_2_io_ipinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_2_io_opinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_2_io_ipinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_2_io_opinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_2_io_ipinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_2_io_ipinSE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_2_io_opinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_2_io_ipinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_2_io_ipinSW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_2_io_opinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_2_io_itrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_2_io_otrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_2_io_itrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_2_io_otrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_2_io_itrackS_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_2_io_otrackS_0; // @[CGRA.scala 273:21]
  wire  gibs_3_clock; // @[CGRA.scala 273:21]
  wire  gibs_3_reset; // @[CGRA.scala 273:21]
  wire  gibs_3_io_cfg_en; // @[CGRA.scala 273:21]
  wire [11:0] gibs_3_io_cfg_addr; // @[CGRA.scala 273:21]
  wire [31:0] gibs_3_io_cfg_data; // @[CGRA.scala 273:21]
  wire [31:0] gibs_3_io_ipinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_3_io_opinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_3_io_ipinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_3_io_opinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_3_io_ipinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_3_io_ipinSE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_3_io_opinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_3_io_ipinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_3_io_ipinSW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_3_io_opinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_3_io_itrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_3_io_otrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_3_io_itrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_3_io_otrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_3_io_itrackS_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_3_io_otrackS_0; // @[CGRA.scala 273:21]
  wire  gibs_4_clock; // @[CGRA.scala 273:21]
  wire  gibs_4_reset; // @[CGRA.scala 273:21]
  wire  gibs_4_io_cfg_en; // @[CGRA.scala 273:21]
  wire [11:0] gibs_4_io_cfg_addr; // @[CGRA.scala 273:21]
  wire [31:0] gibs_4_io_cfg_data; // @[CGRA.scala 273:21]
  wire [31:0] gibs_4_io_ipinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_4_io_opinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_4_io_ipinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_4_io_opinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_4_io_ipinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_4_io_ipinSE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_4_io_opinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_4_io_ipinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_4_io_ipinSW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_4_io_opinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_4_io_itrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_4_io_otrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_4_io_itrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_4_io_otrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_4_io_itrackS_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_4_io_otrackS_0; // @[CGRA.scala 273:21]
  wire  gibs_5_clock; // @[CGRA.scala 273:21]
  wire  gibs_5_reset; // @[CGRA.scala 273:21]
  wire  gibs_5_io_cfg_en; // @[CGRA.scala 273:21]
  wire [11:0] gibs_5_io_cfg_addr; // @[CGRA.scala 273:21]
  wire [31:0] gibs_5_io_cfg_data; // @[CGRA.scala 273:21]
  wire [31:0] gibs_5_io_ipinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_5_io_opinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_5_io_ipinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_5_io_opinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_5_io_ipinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_5_io_ipinSE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_5_io_opinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_5_io_ipinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_5_io_ipinSW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_5_io_opinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_5_io_itrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_5_io_otrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_5_io_itrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_5_io_otrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_5_io_itrackS_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_5_io_otrackS_0; // @[CGRA.scala 273:21]
  wire  gibs_6_clock; // @[CGRA.scala 273:21]
  wire  gibs_6_reset; // @[CGRA.scala 273:21]
  wire  gibs_6_io_cfg_en; // @[CGRA.scala 273:21]
  wire [11:0] gibs_6_io_cfg_addr; // @[CGRA.scala 273:21]
  wire [31:0] gibs_6_io_cfg_data; // @[CGRA.scala 273:21]
  wire [31:0] gibs_6_io_ipinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_6_io_opinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_6_io_ipinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_6_io_opinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_6_io_ipinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_6_io_ipinSE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_6_io_opinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_6_io_ipinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_6_io_ipinSW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_6_io_opinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_6_io_itrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_6_io_otrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_6_io_itrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_6_io_otrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_6_io_itrackS_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_6_io_otrackS_0; // @[CGRA.scala 273:21]
  wire  gibs_7_clock; // @[CGRA.scala 273:21]
  wire  gibs_7_reset; // @[CGRA.scala 273:21]
  wire  gibs_7_io_cfg_en; // @[CGRA.scala 273:21]
  wire [11:0] gibs_7_io_cfg_addr; // @[CGRA.scala 273:21]
  wire [31:0] gibs_7_io_cfg_data; // @[CGRA.scala 273:21]
  wire [31:0] gibs_7_io_ipinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_7_io_opinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_7_io_ipinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_7_io_opinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_7_io_ipinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_7_io_ipinSE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_7_io_opinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_7_io_ipinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_7_io_ipinSW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_7_io_opinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_7_io_itrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_7_io_otrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_7_io_itrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_7_io_otrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_7_io_itrackS_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_7_io_otrackS_0; // @[CGRA.scala 273:21]
  wire  gibs_8_clock; // @[CGRA.scala 273:21]
  wire  gibs_8_reset; // @[CGRA.scala 273:21]
  wire  gibs_8_io_cfg_en; // @[CGRA.scala 273:21]
  wire [11:0] gibs_8_io_cfg_addr; // @[CGRA.scala 273:21]
  wire [31:0] gibs_8_io_cfg_data; // @[CGRA.scala 273:21]
  wire [31:0] gibs_8_io_ipinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_8_io_opinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_8_io_ipinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_8_io_ipinSW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_8_io_opinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_8_io_itrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_8_io_otrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_8_io_itrackS_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_8_io_otrackS_0; // @[CGRA.scala 273:21]
  wire  gibs_9_clock; // @[CGRA.scala 273:21]
  wire  gibs_9_reset; // @[CGRA.scala 273:21]
  wire  gibs_9_io_cfg_en; // @[CGRA.scala 273:21]
  wire [11:0] gibs_9_io_cfg_addr; // @[CGRA.scala 273:21]
  wire [31:0] gibs_9_io_cfg_data; // @[CGRA.scala 273:21]
  wire [31:0] gibs_9_io_ipinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_9_io_ipinNE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_9_io_opinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_9_io_ipinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_9_io_ipinSE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_9_io_opinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_9_io_itrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_9_io_otrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_9_io_itrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_9_io_otrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_9_io_itrackS_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_9_io_otrackS_0; // @[CGRA.scala 273:21]
  wire  gibs_10_clock; // @[CGRA.scala 273:21]
  wire  gibs_10_reset; // @[CGRA.scala 273:21]
  wire  gibs_10_io_cfg_en; // @[CGRA.scala 273:21]
  wire [11:0] gibs_10_io_cfg_addr; // @[CGRA.scala 273:21]
  wire [31:0] gibs_10_io_cfg_data; // @[CGRA.scala 273:21]
  wire [31:0] gibs_10_io_ipinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_10_io_ipinNW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_10_io_opinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_10_io_ipinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_10_io_ipinNE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_10_io_opinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_10_io_ipinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_10_io_ipinSE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_10_io_opinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_10_io_ipinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_10_io_ipinSW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_10_io_opinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_10_io_itrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_10_io_otrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_10_io_itrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_10_io_otrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_10_io_itrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_10_io_otrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_10_io_itrackS_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_10_io_otrackS_0; // @[CGRA.scala 273:21]
  wire  gibs_11_clock; // @[CGRA.scala 273:21]
  wire  gibs_11_reset; // @[CGRA.scala 273:21]
  wire  gibs_11_io_cfg_en; // @[CGRA.scala 273:21]
  wire [11:0] gibs_11_io_cfg_addr; // @[CGRA.scala 273:21]
  wire [31:0] gibs_11_io_cfg_data; // @[CGRA.scala 273:21]
  wire [31:0] gibs_11_io_ipinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_11_io_ipinNW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_11_io_opinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_11_io_ipinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_11_io_ipinNE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_11_io_opinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_11_io_ipinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_11_io_ipinSE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_11_io_opinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_11_io_ipinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_11_io_ipinSW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_11_io_opinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_11_io_itrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_11_io_otrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_11_io_itrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_11_io_otrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_11_io_itrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_11_io_otrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_11_io_itrackS_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_11_io_otrackS_0; // @[CGRA.scala 273:21]
  wire  gibs_12_clock; // @[CGRA.scala 273:21]
  wire  gibs_12_reset; // @[CGRA.scala 273:21]
  wire  gibs_12_io_cfg_en; // @[CGRA.scala 273:21]
  wire [11:0] gibs_12_io_cfg_addr; // @[CGRA.scala 273:21]
  wire [31:0] gibs_12_io_cfg_data; // @[CGRA.scala 273:21]
  wire [31:0] gibs_12_io_ipinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_12_io_ipinNW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_12_io_opinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_12_io_ipinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_12_io_ipinNE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_12_io_opinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_12_io_ipinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_12_io_ipinSE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_12_io_opinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_12_io_ipinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_12_io_ipinSW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_12_io_opinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_12_io_itrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_12_io_otrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_12_io_itrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_12_io_otrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_12_io_itrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_12_io_otrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_12_io_itrackS_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_12_io_otrackS_0; // @[CGRA.scala 273:21]
  wire  gibs_13_clock; // @[CGRA.scala 273:21]
  wire  gibs_13_reset; // @[CGRA.scala 273:21]
  wire  gibs_13_io_cfg_en; // @[CGRA.scala 273:21]
  wire [11:0] gibs_13_io_cfg_addr; // @[CGRA.scala 273:21]
  wire [31:0] gibs_13_io_cfg_data; // @[CGRA.scala 273:21]
  wire [31:0] gibs_13_io_ipinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_13_io_ipinNW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_13_io_opinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_13_io_ipinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_13_io_ipinNE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_13_io_opinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_13_io_ipinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_13_io_ipinSE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_13_io_opinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_13_io_ipinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_13_io_ipinSW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_13_io_opinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_13_io_itrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_13_io_otrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_13_io_itrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_13_io_otrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_13_io_itrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_13_io_otrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_13_io_itrackS_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_13_io_otrackS_0; // @[CGRA.scala 273:21]
  wire  gibs_14_clock; // @[CGRA.scala 273:21]
  wire  gibs_14_reset; // @[CGRA.scala 273:21]
  wire  gibs_14_io_cfg_en; // @[CGRA.scala 273:21]
  wire [11:0] gibs_14_io_cfg_addr; // @[CGRA.scala 273:21]
  wire [31:0] gibs_14_io_cfg_data; // @[CGRA.scala 273:21]
  wire [31:0] gibs_14_io_ipinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_14_io_ipinNW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_14_io_opinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_14_io_ipinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_14_io_ipinNE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_14_io_opinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_14_io_ipinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_14_io_ipinSE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_14_io_opinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_14_io_ipinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_14_io_ipinSW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_14_io_opinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_14_io_itrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_14_io_otrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_14_io_itrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_14_io_otrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_14_io_itrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_14_io_otrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_14_io_itrackS_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_14_io_otrackS_0; // @[CGRA.scala 273:21]
  wire  gibs_15_clock; // @[CGRA.scala 273:21]
  wire  gibs_15_reset; // @[CGRA.scala 273:21]
  wire  gibs_15_io_cfg_en; // @[CGRA.scala 273:21]
  wire [11:0] gibs_15_io_cfg_addr; // @[CGRA.scala 273:21]
  wire [31:0] gibs_15_io_cfg_data; // @[CGRA.scala 273:21]
  wire [31:0] gibs_15_io_ipinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_15_io_ipinNW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_15_io_opinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_15_io_ipinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_15_io_ipinNE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_15_io_opinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_15_io_ipinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_15_io_ipinSE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_15_io_opinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_15_io_ipinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_15_io_ipinSW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_15_io_opinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_15_io_itrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_15_io_otrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_15_io_itrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_15_io_otrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_15_io_itrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_15_io_otrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_15_io_itrackS_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_15_io_otrackS_0; // @[CGRA.scala 273:21]
  wire  gibs_16_clock; // @[CGRA.scala 273:21]
  wire  gibs_16_reset; // @[CGRA.scala 273:21]
  wire  gibs_16_io_cfg_en; // @[CGRA.scala 273:21]
  wire [11:0] gibs_16_io_cfg_addr; // @[CGRA.scala 273:21]
  wire [31:0] gibs_16_io_cfg_data; // @[CGRA.scala 273:21]
  wire [31:0] gibs_16_io_ipinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_16_io_ipinNW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_16_io_opinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_16_io_ipinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_16_io_ipinNE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_16_io_opinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_16_io_ipinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_16_io_ipinSE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_16_io_opinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_16_io_ipinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_16_io_ipinSW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_16_io_opinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_16_io_itrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_16_io_otrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_16_io_itrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_16_io_otrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_16_io_itrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_16_io_otrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_16_io_itrackS_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_16_io_otrackS_0; // @[CGRA.scala 273:21]
  wire  gibs_17_clock; // @[CGRA.scala 273:21]
  wire  gibs_17_reset; // @[CGRA.scala 273:21]
  wire  gibs_17_io_cfg_en; // @[CGRA.scala 273:21]
  wire [11:0] gibs_17_io_cfg_addr; // @[CGRA.scala 273:21]
  wire [31:0] gibs_17_io_cfg_data; // @[CGRA.scala 273:21]
  wire [31:0] gibs_17_io_ipinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_17_io_ipinNW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_17_io_opinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_17_io_ipinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_17_io_ipinSW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_17_io_opinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_17_io_itrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_17_io_otrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_17_io_itrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_17_io_otrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_17_io_itrackS_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_17_io_otrackS_0; // @[CGRA.scala 273:21]
  wire  gibs_18_clock; // @[CGRA.scala 273:21]
  wire  gibs_18_reset; // @[CGRA.scala 273:21]
  wire  gibs_18_io_cfg_en; // @[CGRA.scala 273:21]
  wire [11:0] gibs_18_io_cfg_addr; // @[CGRA.scala 273:21]
  wire [31:0] gibs_18_io_cfg_data; // @[CGRA.scala 273:21]
  wire [31:0] gibs_18_io_ipinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_18_io_ipinNE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_18_io_opinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_18_io_ipinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_18_io_ipinSE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_18_io_opinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_18_io_itrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_18_io_otrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_18_io_itrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_18_io_otrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_18_io_itrackS_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_18_io_otrackS_0; // @[CGRA.scala 273:21]
  wire  gibs_19_clock; // @[CGRA.scala 273:21]
  wire  gibs_19_reset; // @[CGRA.scala 273:21]
  wire  gibs_19_io_cfg_en; // @[CGRA.scala 273:21]
  wire [11:0] gibs_19_io_cfg_addr; // @[CGRA.scala 273:21]
  wire [31:0] gibs_19_io_cfg_data; // @[CGRA.scala 273:21]
  wire [31:0] gibs_19_io_ipinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_19_io_ipinNW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_19_io_opinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_19_io_ipinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_19_io_ipinNE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_19_io_opinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_19_io_ipinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_19_io_ipinSE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_19_io_opinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_19_io_ipinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_19_io_ipinSW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_19_io_opinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_19_io_itrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_19_io_otrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_19_io_itrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_19_io_otrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_19_io_itrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_19_io_otrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_19_io_itrackS_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_19_io_otrackS_0; // @[CGRA.scala 273:21]
  wire  gibs_20_clock; // @[CGRA.scala 273:21]
  wire  gibs_20_reset; // @[CGRA.scala 273:21]
  wire  gibs_20_io_cfg_en; // @[CGRA.scala 273:21]
  wire [11:0] gibs_20_io_cfg_addr; // @[CGRA.scala 273:21]
  wire [31:0] gibs_20_io_cfg_data; // @[CGRA.scala 273:21]
  wire [31:0] gibs_20_io_ipinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_20_io_ipinNW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_20_io_opinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_20_io_ipinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_20_io_ipinNE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_20_io_opinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_20_io_ipinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_20_io_ipinSE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_20_io_opinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_20_io_ipinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_20_io_ipinSW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_20_io_opinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_20_io_itrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_20_io_otrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_20_io_itrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_20_io_otrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_20_io_itrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_20_io_otrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_20_io_itrackS_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_20_io_otrackS_0; // @[CGRA.scala 273:21]
  wire  gibs_21_clock; // @[CGRA.scala 273:21]
  wire  gibs_21_reset; // @[CGRA.scala 273:21]
  wire  gibs_21_io_cfg_en; // @[CGRA.scala 273:21]
  wire [11:0] gibs_21_io_cfg_addr; // @[CGRA.scala 273:21]
  wire [31:0] gibs_21_io_cfg_data; // @[CGRA.scala 273:21]
  wire [31:0] gibs_21_io_ipinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_21_io_ipinNW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_21_io_opinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_21_io_ipinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_21_io_ipinNE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_21_io_opinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_21_io_ipinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_21_io_ipinSE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_21_io_opinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_21_io_ipinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_21_io_ipinSW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_21_io_opinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_21_io_itrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_21_io_otrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_21_io_itrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_21_io_otrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_21_io_itrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_21_io_otrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_21_io_itrackS_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_21_io_otrackS_0; // @[CGRA.scala 273:21]
  wire  gibs_22_clock; // @[CGRA.scala 273:21]
  wire  gibs_22_reset; // @[CGRA.scala 273:21]
  wire  gibs_22_io_cfg_en; // @[CGRA.scala 273:21]
  wire [11:0] gibs_22_io_cfg_addr; // @[CGRA.scala 273:21]
  wire [31:0] gibs_22_io_cfg_data; // @[CGRA.scala 273:21]
  wire [31:0] gibs_22_io_ipinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_22_io_ipinNW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_22_io_opinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_22_io_ipinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_22_io_ipinNE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_22_io_opinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_22_io_ipinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_22_io_ipinSE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_22_io_opinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_22_io_ipinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_22_io_ipinSW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_22_io_opinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_22_io_itrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_22_io_otrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_22_io_itrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_22_io_otrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_22_io_itrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_22_io_otrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_22_io_itrackS_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_22_io_otrackS_0; // @[CGRA.scala 273:21]
  wire  gibs_23_clock; // @[CGRA.scala 273:21]
  wire  gibs_23_reset; // @[CGRA.scala 273:21]
  wire  gibs_23_io_cfg_en; // @[CGRA.scala 273:21]
  wire [11:0] gibs_23_io_cfg_addr; // @[CGRA.scala 273:21]
  wire [31:0] gibs_23_io_cfg_data; // @[CGRA.scala 273:21]
  wire [31:0] gibs_23_io_ipinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_23_io_ipinNW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_23_io_opinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_23_io_ipinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_23_io_ipinNE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_23_io_opinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_23_io_ipinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_23_io_ipinSE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_23_io_opinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_23_io_ipinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_23_io_ipinSW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_23_io_opinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_23_io_itrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_23_io_otrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_23_io_itrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_23_io_otrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_23_io_itrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_23_io_otrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_23_io_itrackS_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_23_io_otrackS_0; // @[CGRA.scala 273:21]
  wire  gibs_24_clock; // @[CGRA.scala 273:21]
  wire  gibs_24_reset; // @[CGRA.scala 273:21]
  wire  gibs_24_io_cfg_en; // @[CGRA.scala 273:21]
  wire [11:0] gibs_24_io_cfg_addr; // @[CGRA.scala 273:21]
  wire [31:0] gibs_24_io_cfg_data; // @[CGRA.scala 273:21]
  wire [31:0] gibs_24_io_ipinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_24_io_ipinNW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_24_io_opinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_24_io_ipinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_24_io_ipinNE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_24_io_opinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_24_io_ipinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_24_io_ipinSE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_24_io_opinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_24_io_ipinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_24_io_ipinSW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_24_io_opinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_24_io_itrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_24_io_otrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_24_io_itrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_24_io_otrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_24_io_itrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_24_io_otrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_24_io_itrackS_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_24_io_otrackS_0; // @[CGRA.scala 273:21]
  wire  gibs_25_clock; // @[CGRA.scala 273:21]
  wire  gibs_25_reset; // @[CGRA.scala 273:21]
  wire  gibs_25_io_cfg_en; // @[CGRA.scala 273:21]
  wire [11:0] gibs_25_io_cfg_addr; // @[CGRA.scala 273:21]
  wire [31:0] gibs_25_io_cfg_data; // @[CGRA.scala 273:21]
  wire [31:0] gibs_25_io_ipinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_25_io_ipinNW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_25_io_opinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_25_io_ipinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_25_io_ipinNE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_25_io_opinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_25_io_ipinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_25_io_ipinSE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_25_io_opinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_25_io_ipinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_25_io_ipinSW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_25_io_opinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_25_io_itrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_25_io_otrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_25_io_itrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_25_io_otrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_25_io_itrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_25_io_otrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_25_io_itrackS_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_25_io_otrackS_0; // @[CGRA.scala 273:21]
  wire  gibs_26_clock; // @[CGRA.scala 273:21]
  wire  gibs_26_reset; // @[CGRA.scala 273:21]
  wire  gibs_26_io_cfg_en; // @[CGRA.scala 273:21]
  wire [11:0] gibs_26_io_cfg_addr; // @[CGRA.scala 273:21]
  wire [31:0] gibs_26_io_cfg_data; // @[CGRA.scala 273:21]
  wire [31:0] gibs_26_io_ipinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_26_io_ipinNW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_26_io_opinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_26_io_ipinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_26_io_ipinSW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_26_io_opinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_26_io_itrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_26_io_otrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_26_io_itrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_26_io_otrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_26_io_itrackS_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_26_io_otrackS_0; // @[CGRA.scala 273:21]
  wire  gibs_27_clock; // @[CGRA.scala 273:21]
  wire  gibs_27_reset; // @[CGRA.scala 273:21]
  wire  gibs_27_io_cfg_en; // @[CGRA.scala 273:21]
  wire [11:0] gibs_27_io_cfg_addr; // @[CGRA.scala 273:21]
  wire [31:0] gibs_27_io_cfg_data; // @[CGRA.scala 273:21]
  wire [31:0] gibs_27_io_ipinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_27_io_ipinNE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_27_io_opinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_27_io_ipinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_27_io_ipinSE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_27_io_opinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_27_io_itrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_27_io_otrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_27_io_itrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_27_io_otrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_27_io_itrackS_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_27_io_otrackS_0; // @[CGRA.scala 273:21]
  wire  gibs_28_clock; // @[CGRA.scala 273:21]
  wire  gibs_28_reset; // @[CGRA.scala 273:21]
  wire  gibs_28_io_cfg_en; // @[CGRA.scala 273:21]
  wire [11:0] gibs_28_io_cfg_addr; // @[CGRA.scala 273:21]
  wire [31:0] gibs_28_io_cfg_data; // @[CGRA.scala 273:21]
  wire [31:0] gibs_28_io_ipinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_28_io_ipinNW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_28_io_opinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_28_io_ipinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_28_io_ipinNE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_28_io_opinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_28_io_ipinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_28_io_ipinSE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_28_io_opinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_28_io_ipinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_28_io_ipinSW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_28_io_opinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_28_io_itrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_28_io_otrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_28_io_itrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_28_io_otrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_28_io_itrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_28_io_otrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_28_io_itrackS_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_28_io_otrackS_0; // @[CGRA.scala 273:21]
  wire  gibs_29_clock; // @[CGRA.scala 273:21]
  wire  gibs_29_reset; // @[CGRA.scala 273:21]
  wire  gibs_29_io_cfg_en; // @[CGRA.scala 273:21]
  wire [11:0] gibs_29_io_cfg_addr; // @[CGRA.scala 273:21]
  wire [31:0] gibs_29_io_cfg_data; // @[CGRA.scala 273:21]
  wire [31:0] gibs_29_io_ipinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_29_io_ipinNW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_29_io_opinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_29_io_ipinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_29_io_ipinNE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_29_io_opinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_29_io_ipinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_29_io_ipinSE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_29_io_opinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_29_io_ipinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_29_io_ipinSW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_29_io_opinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_29_io_itrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_29_io_otrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_29_io_itrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_29_io_otrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_29_io_itrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_29_io_otrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_29_io_itrackS_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_29_io_otrackS_0; // @[CGRA.scala 273:21]
  wire  gibs_30_clock; // @[CGRA.scala 273:21]
  wire  gibs_30_reset; // @[CGRA.scala 273:21]
  wire  gibs_30_io_cfg_en; // @[CGRA.scala 273:21]
  wire [11:0] gibs_30_io_cfg_addr; // @[CGRA.scala 273:21]
  wire [31:0] gibs_30_io_cfg_data; // @[CGRA.scala 273:21]
  wire [31:0] gibs_30_io_ipinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_30_io_ipinNW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_30_io_opinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_30_io_ipinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_30_io_ipinNE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_30_io_opinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_30_io_ipinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_30_io_ipinSE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_30_io_opinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_30_io_ipinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_30_io_ipinSW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_30_io_opinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_30_io_itrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_30_io_otrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_30_io_itrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_30_io_otrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_30_io_itrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_30_io_otrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_30_io_itrackS_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_30_io_otrackS_0; // @[CGRA.scala 273:21]
  wire  gibs_31_clock; // @[CGRA.scala 273:21]
  wire  gibs_31_reset; // @[CGRA.scala 273:21]
  wire  gibs_31_io_cfg_en; // @[CGRA.scala 273:21]
  wire [11:0] gibs_31_io_cfg_addr; // @[CGRA.scala 273:21]
  wire [31:0] gibs_31_io_cfg_data; // @[CGRA.scala 273:21]
  wire [31:0] gibs_31_io_ipinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_31_io_ipinNW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_31_io_opinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_31_io_ipinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_31_io_ipinNE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_31_io_opinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_31_io_ipinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_31_io_ipinSE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_31_io_opinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_31_io_ipinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_31_io_ipinSW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_31_io_opinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_31_io_itrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_31_io_otrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_31_io_itrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_31_io_otrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_31_io_itrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_31_io_otrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_31_io_itrackS_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_31_io_otrackS_0; // @[CGRA.scala 273:21]
  wire  gibs_32_clock; // @[CGRA.scala 273:21]
  wire  gibs_32_reset; // @[CGRA.scala 273:21]
  wire  gibs_32_io_cfg_en; // @[CGRA.scala 273:21]
  wire [11:0] gibs_32_io_cfg_addr; // @[CGRA.scala 273:21]
  wire [31:0] gibs_32_io_cfg_data; // @[CGRA.scala 273:21]
  wire [31:0] gibs_32_io_ipinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_32_io_ipinNW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_32_io_opinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_32_io_ipinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_32_io_ipinNE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_32_io_opinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_32_io_ipinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_32_io_ipinSE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_32_io_opinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_32_io_ipinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_32_io_ipinSW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_32_io_opinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_32_io_itrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_32_io_otrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_32_io_itrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_32_io_otrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_32_io_itrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_32_io_otrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_32_io_itrackS_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_32_io_otrackS_0; // @[CGRA.scala 273:21]
  wire  gibs_33_clock; // @[CGRA.scala 273:21]
  wire  gibs_33_reset; // @[CGRA.scala 273:21]
  wire  gibs_33_io_cfg_en; // @[CGRA.scala 273:21]
  wire [11:0] gibs_33_io_cfg_addr; // @[CGRA.scala 273:21]
  wire [31:0] gibs_33_io_cfg_data; // @[CGRA.scala 273:21]
  wire [31:0] gibs_33_io_ipinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_33_io_ipinNW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_33_io_opinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_33_io_ipinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_33_io_ipinNE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_33_io_opinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_33_io_ipinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_33_io_ipinSE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_33_io_opinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_33_io_ipinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_33_io_ipinSW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_33_io_opinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_33_io_itrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_33_io_otrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_33_io_itrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_33_io_otrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_33_io_itrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_33_io_otrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_33_io_itrackS_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_33_io_otrackS_0; // @[CGRA.scala 273:21]
  wire  gibs_34_clock; // @[CGRA.scala 273:21]
  wire  gibs_34_reset; // @[CGRA.scala 273:21]
  wire  gibs_34_io_cfg_en; // @[CGRA.scala 273:21]
  wire [11:0] gibs_34_io_cfg_addr; // @[CGRA.scala 273:21]
  wire [31:0] gibs_34_io_cfg_data; // @[CGRA.scala 273:21]
  wire [31:0] gibs_34_io_ipinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_34_io_ipinNW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_34_io_opinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_34_io_ipinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_34_io_ipinNE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_34_io_opinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_34_io_ipinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_34_io_ipinSE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_34_io_opinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_34_io_ipinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_34_io_ipinSW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_34_io_opinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_34_io_itrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_34_io_otrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_34_io_itrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_34_io_otrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_34_io_itrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_34_io_otrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_34_io_itrackS_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_34_io_otrackS_0; // @[CGRA.scala 273:21]
  wire  gibs_35_clock; // @[CGRA.scala 273:21]
  wire  gibs_35_reset; // @[CGRA.scala 273:21]
  wire  gibs_35_io_cfg_en; // @[CGRA.scala 273:21]
  wire [11:0] gibs_35_io_cfg_addr; // @[CGRA.scala 273:21]
  wire [31:0] gibs_35_io_cfg_data; // @[CGRA.scala 273:21]
  wire [31:0] gibs_35_io_ipinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_35_io_ipinNW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_35_io_opinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_35_io_ipinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_35_io_ipinSW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_35_io_opinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_35_io_itrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_35_io_otrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_35_io_itrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_35_io_otrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_35_io_itrackS_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_35_io_otrackS_0; // @[CGRA.scala 273:21]
  wire  gibs_36_clock; // @[CGRA.scala 273:21]
  wire  gibs_36_reset; // @[CGRA.scala 273:21]
  wire  gibs_36_io_cfg_en; // @[CGRA.scala 273:21]
  wire [11:0] gibs_36_io_cfg_addr; // @[CGRA.scala 273:21]
  wire [31:0] gibs_36_io_cfg_data; // @[CGRA.scala 273:21]
  wire [31:0] gibs_36_io_ipinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_36_io_ipinNE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_36_io_opinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_36_io_ipinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_36_io_ipinSE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_36_io_opinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_36_io_itrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_36_io_otrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_36_io_itrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_36_io_otrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_36_io_itrackS_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_36_io_otrackS_0; // @[CGRA.scala 273:21]
  wire  gibs_37_clock; // @[CGRA.scala 273:21]
  wire  gibs_37_reset; // @[CGRA.scala 273:21]
  wire  gibs_37_io_cfg_en; // @[CGRA.scala 273:21]
  wire [11:0] gibs_37_io_cfg_addr; // @[CGRA.scala 273:21]
  wire [31:0] gibs_37_io_cfg_data; // @[CGRA.scala 273:21]
  wire [31:0] gibs_37_io_ipinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_37_io_ipinNW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_37_io_opinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_37_io_ipinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_37_io_ipinNE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_37_io_opinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_37_io_ipinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_37_io_ipinSE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_37_io_opinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_37_io_ipinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_37_io_ipinSW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_37_io_opinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_37_io_itrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_37_io_otrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_37_io_itrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_37_io_otrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_37_io_itrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_37_io_otrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_37_io_itrackS_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_37_io_otrackS_0; // @[CGRA.scala 273:21]
  wire  gibs_38_clock; // @[CGRA.scala 273:21]
  wire  gibs_38_reset; // @[CGRA.scala 273:21]
  wire  gibs_38_io_cfg_en; // @[CGRA.scala 273:21]
  wire [11:0] gibs_38_io_cfg_addr; // @[CGRA.scala 273:21]
  wire [31:0] gibs_38_io_cfg_data; // @[CGRA.scala 273:21]
  wire [31:0] gibs_38_io_ipinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_38_io_ipinNW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_38_io_opinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_38_io_ipinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_38_io_ipinNE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_38_io_opinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_38_io_ipinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_38_io_ipinSE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_38_io_opinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_38_io_ipinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_38_io_ipinSW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_38_io_opinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_38_io_itrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_38_io_otrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_38_io_itrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_38_io_otrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_38_io_itrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_38_io_otrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_38_io_itrackS_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_38_io_otrackS_0; // @[CGRA.scala 273:21]
  wire  gibs_39_clock; // @[CGRA.scala 273:21]
  wire  gibs_39_reset; // @[CGRA.scala 273:21]
  wire  gibs_39_io_cfg_en; // @[CGRA.scala 273:21]
  wire [11:0] gibs_39_io_cfg_addr; // @[CGRA.scala 273:21]
  wire [31:0] gibs_39_io_cfg_data; // @[CGRA.scala 273:21]
  wire [31:0] gibs_39_io_ipinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_39_io_ipinNW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_39_io_opinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_39_io_ipinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_39_io_ipinNE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_39_io_opinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_39_io_ipinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_39_io_ipinSE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_39_io_opinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_39_io_ipinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_39_io_ipinSW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_39_io_opinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_39_io_itrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_39_io_otrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_39_io_itrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_39_io_otrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_39_io_itrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_39_io_otrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_39_io_itrackS_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_39_io_otrackS_0; // @[CGRA.scala 273:21]
  wire  gibs_40_clock; // @[CGRA.scala 273:21]
  wire  gibs_40_reset; // @[CGRA.scala 273:21]
  wire  gibs_40_io_cfg_en; // @[CGRA.scala 273:21]
  wire [11:0] gibs_40_io_cfg_addr; // @[CGRA.scala 273:21]
  wire [31:0] gibs_40_io_cfg_data; // @[CGRA.scala 273:21]
  wire [31:0] gibs_40_io_ipinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_40_io_ipinNW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_40_io_opinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_40_io_ipinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_40_io_ipinNE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_40_io_opinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_40_io_ipinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_40_io_ipinSE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_40_io_opinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_40_io_ipinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_40_io_ipinSW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_40_io_opinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_40_io_itrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_40_io_otrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_40_io_itrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_40_io_otrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_40_io_itrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_40_io_otrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_40_io_itrackS_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_40_io_otrackS_0; // @[CGRA.scala 273:21]
  wire  gibs_41_clock; // @[CGRA.scala 273:21]
  wire  gibs_41_reset; // @[CGRA.scala 273:21]
  wire  gibs_41_io_cfg_en; // @[CGRA.scala 273:21]
  wire [11:0] gibs_41_io_cfg_addr; // @[CGRA.scala 273:21]
  wire [31:0] gibs_41_io_cfg_data; // @[CGRA.scala 273:21]
  wire [31:0] gibs_41_io_ipinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_41_io_ipinNW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_41_io_opinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_41_io_ipinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_41_io_ipinNE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_41_io_opinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_41_io_ipinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_41_io_ipinSE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_41_io_opinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_41_io_ipinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_41_io_ipinSW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_41_io_opinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_41_io_itrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_41_io_otrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_41_io_itrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_41_io_otrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_41_io_itrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_41_io_otrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_41_io_itrackS_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_41_io_otrackS_0; // @[CGRA.scala 273:21]
  wire  gibs_42_clock; // @[CGRA.scala 273:21]
  wire  gibs_42_reset; // @[CGRA.scala 273:21]
  wire  gibs_42_io_cfg_en; // @[CGRA.scala 273:21]
  wire [11:0] gibs_42_io_cfg_addr; // @[CGRA.scala 273:21]
  wire [31:0] gibs_42_io_cfg_data; // @[CGRA.scala 273:21]
  wire [31:0] gibs_42_io_ipinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_42_io_ipinNW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_42_io_opinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_42_io_ipinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_42_io_ipinNE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_42_io_opinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_42_io_ipinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_42_io_ipinSE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_42_io_opinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_42_io_ipinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_42_io_ipinSW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_42_io_opinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_42_io_itrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_42_io_otrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_42_io_itrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_42_io_otrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_42_io_itrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_42_io_otrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_42_io_itrackS_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_42_io_otrackS_0; // @[CGRA.scala 273:21]
  wire  gibs_43_clock; // @[CGRA.scala 273:21]
  wire  gibs_43_reset; // @[CGRA.scala 273:21]
  wire  gibs_43_io_cfg_en; // @[CGRA.scala 273:21]
  wire [11:0] gibs_43_io_cfg_addr; // @[CGRA.scala 273:21]
  wire [31:0] gibs_43_io_cfg_data; // @[CGRA.scala 273:21]
  wire [31:0] gibs_43_io_ipinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_43_io_ipinNW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_43_io_opinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_43_io_ipinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_43_io_ipinNE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_43_io_opinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_43_io_ipinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_43_io_ipinSE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_43_io_opinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_43_io_ipinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_43_io_ipinSW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_43_io_opinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_43_io_itrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_43_io_otrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_43_io_itrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_43_io_otrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_43_io_itrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_43_io_otrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_43_io_itrackS_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_43_io_otrackS_0; // @[CGRA.scala 273:21]
  wire  gibs_44_clock; // @[CGRA.scala 273:21]
  wire  gibs_44_reset; // @[CGRA.scala 273:21]
  wire  gibs_44_io_cfg_en; // @[CGRA.scala 273:21]
  wire [11:0] gibs_44_io_cfg_addr; // @[CGRA.scala 273:21]
  wire [31:0] gibs_44_io_cfg_data; // @[CGRA.scala 273:21]
  wire [31:0] gibs_44_io_ipinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_44_io_ipinNW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_44_io_opinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_44_io_ipinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_44_io_ipinSW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_44_io_opinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_44_io_itrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_44_io_otrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_44_io_itrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_44_io_otrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_44_io_itrackS_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_44_io_otrackS_0; // @[CGRA.scala 273:21]
  wire  gibs_45_clock; // @[CGRA.scala 273:21]
  wire  gibs_45_reset; // @[CGRA.scala 273:21]
  wire  gibs_45_io_cfg_en; // @[CGRA.scala 273:21]
  wire [11:0] gibs_45_io_cfg_addr; // @[CGRA.scala 273:21]
  wire [31:0] gibs_45_io_cfg_data; // @[CGRA.scala 273:21]
  wire [31:0] gibs_45_io_ipinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_45_io_ipinNE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_45_io_opinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_45_io_ipinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_45_io_ipinSE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_45_io_opinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_45_io_itrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_45_io_otrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_45_io_itrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_45_io_otrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_45_io_itrackS_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_45_io_otrackS_0; // @[CGRA.scala 273:21]
  wire  gibs_46_clock; // @[CGRA.scala 273:21]
  wire  gibs_46_reset; // @[CGRA.scala 273:21]
  wire  gibs_46_io_cfg_en; // @[CGRA.scala 273:21]
  wire [11:0] gibs_46_io_cfg_addr; // @[CGRA.scala 273:21]
  wire [31:0] gibs_46_io_cfg_data; // @[CGRA.scala 273:21]
  wire [31:0] gibs_46_io_ipinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_46_io_ipinNW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_46_io_opinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_46_io_ipinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_46_io_ipinNE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_46_io_opinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_46_io_ipinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_46_io_ipinSE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_46_io_opinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_46_io_ipinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_46_io_ipinSW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_46_io_opinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_46_io_itrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_46_io_otrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_46_io_itrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_46_io_otrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_46_io_itrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_46_io_otrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_46_io_itrackS_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_46_io_otrackS_0; // @[CGRA.scala 273:21]
  wire  gibs_47_clock; // @[CGRA.scala 273:21]
  wire  gibs_47_reset; // @[CGRA.scala 273:21]
  wire  gibs_47_io_cfg_en; // @[CGRA.scala 273:21]
  wire [11:0] gibs_47_io_cfg_addr; // @[CGRA.scala 273:21]
  wire [31:0] gibs_47_io_cfg_data; // @[CGRA.scala 273:21]
  wire [31:0] gibs_47_io_ipinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_47_io_ipinNW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_47_io_opinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_47_io_ipinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_47_io_ipinNE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_47_io_opinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_47_io_ipinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_47_io_ipinSE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_47_io_opinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_47_io_ipinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_47_io_ipinSW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_47_io_opinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_47_io_itrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_47_io_otrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_47_io_itrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_47_io_otrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_47_io_itrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_47_io_otrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_47_io_itrackS_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_47_io_otrackS_0; // @[CGRA.scala 273:21]
  wire  gibs_48_clock; // @[CGRA.scala 273:21]
  wire  gibs_48_reset; // @[CGRA.scala 273:21]
  wire  gibs_48_io_cfg_en; // @[CGRA.scala 273:21]
  wire [11:0] gibs_48_io_cfg_addr; // @[CGRA.scala 273:21]
  wire [31:0] gibs_48_io_cfg_data; // @[CGRA.scala 273:21]
  wire [31:0] gibs_48_io_ipinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_48_io_ipinNW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_48_io_opinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_48_io_ipinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_48_io_ipinNE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_48_io_opinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_48_io_ipinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_48_io_ipinSE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_48_io_opinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_48_io_ipinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_48_io_ipinSW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_48_io_opinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_48_io_itrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_48_io_otrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_48_io_itrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_48_io_otrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_48_io_itrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_48_io_otrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_48_io_itrackS_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_48_io_otrackS_0; // @[CGRA.scala 273:21]
  wire  gibs_49_clock; // @[CGRA.scala 273:21]
  wire  gibs_49_reset; // @[CGRA.scala 273:21]
  wire  gibs_49_io_cfg_en; // @[CGRA.scala 273:21]
  wire [11:0] gibs_49_io_cfg_addr; // @[CGRA.scala 273:21]
  wire [31:0] gibs_49_io_cfg_data; // @[CGRA.scala 273:21]
  wire [31:0] gibs_49_io_ipinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_49_io_ipinNW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_49_io_opinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_49_io_ipinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_49_io_ipinNE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_49_io_opinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_49_io_ipinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_49_io_ipinSE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_49_io_opinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_49_io_ipinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_49_io_ipinSW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_49_io_opinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_49_io_itrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_49_io_otrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_49_io_itrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_49_io_otrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_49_io_itrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_49_io_otrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_49_io_itrackS_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_49_io_otrackS_0; // @[CGRA.scala 273:21]
  wire  gibs_50_clock; // @[CGRA.scala 273:21]
  wire  gibs_50_reset; // @[CGRA.scala 273:21]
  wire  gibs_50_io_cfg_en; // @[CGRA.scala 273:21]
  wire [11:0] gibs_50_io_cfg_addr; // @[CGRA.scala 273:21]
  wire [31:0] gibs_50_io_cfg_data; // @[CGRA.scala 273:21]
  wire [31:0] gibs_50_io_ipinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_50_io_ipinNW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_50_io_opinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_50_io_ipinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_50_io_ipinNE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_50_io_opinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_50_io_ipinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_50_io_ipinSE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_50_io_opinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_50_io_ipinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_50_io_ipinSW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_50_io_opinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_50_io_itrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_50_io_otrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_50_io_itrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_50_io_otrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_50_io_itrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_50_io_otrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_50_io_itrackS_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_50_io_otrackS_0; // @[CGRA.scala 273:21]
  wire  gibs_51_clock; // @[CGRA.scala 273:21]
  wire  gibs_51_reset; // @[CGRA.scala 273:21]
  wire  gibs_51_io_cfg_en; // @[CGRA.scala 273:21]
  wire [11:0] gibs_51_io_cfg_addr; // @[CGRA.scala 273:21]
  wire [31:0] gibs_51_io_cfg_data; // @[CGRA.scala 273:21]
  wire [31:0] gibs_51_io_ipinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_51_io_ipinNW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_51_io_opinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_51_io_ipinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_51_io_ipinNE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_51_io_opinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_51_io_ipinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_51_io_ipinSE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_51_io_opinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_51_io_ipinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_51_io_ipinSW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_51_io_opinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_51_io_itrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_51_io_otrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_51_io_itrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_51_io_otrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_51_io_itrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_51_io_otrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_51_io_itrackS_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_51_io_otrackS_0; // @[CGRA.scala 273:21]
  wire  gibs_52_clock; // @[CGRA.scala 273:21]
  wire  gibs_52_reset; // @[CGRA.scala 273:21]
  wire  gibs_52_io_cfg_en; // @[CGRA.scala 273:21]
  wire [11:0] gibs_52_io_cfg_addr; // @[CGRA.scala 273:21]
  wire [31:0] gibs_52_io_cfg_data; // @[CGRA.scala 273:21]
  wire [31:0] gibs_52_io_ipinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_52_io_ipinNW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_52_io_opinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_52_io_ipinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_52_io_ipinNE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_52_io_opinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_52_io_ipinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_52_io_ipinSE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_52_io_opinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_52_io_ipinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_52_io_ipinSW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_52_io_opinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_52_io_itrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_52_io_otrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_52_io_itrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_52_io_otrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_52_io_itrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_52_io_otrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_52_io_itrackS_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_52_io_otrackS_0; // @[CGRA.scala 273:21]
  wire  gibs_53_clock; // @[CGRA.scala 273:21]
  wire  gibs_53_reset; // @[CGRA.scala 273:21]
  wire  gibs_53_io_cfg_en; // @[CGRA.scala 273:21]
  wire [11:0] gibs_53_io_cfg_addr; // @[CGRA.scala 273:21]
  wire [31:0] gibs_53_io_cfg_data; // @[CGRA.scala 273:21]
  wire [31:0] gibs_53_io_ipinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_53_io_ipinNW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_53_io_opinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_53_io_ipinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_53_io_ipinSW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_53_io_opinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_53_io_itrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_53_io_otrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_53_io_itrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_53_io_otrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_53_io_itrackS_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_53_io_otrackS_0; // @[CGRA.scala 273:21]
  wire  gibs_54_clock; // @[CGRA.scala 273:21]
  wire  gibs_54_reset; // @[CGRA.scala 273:21]
  wire  gibs_54_io_cfg_en; // @[CGRA.scala 273:21]
  wire [11:0] gibs_54_io_cfg_addr; // @[CGRA.scala 273:21]
  wire [31:0] gibs_54_io_cfg_data; // @[CGRA.scala 273:21]
  wire [31:0] gibs_54_io_ipinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_54_io_ipinNE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_54_io_opinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_54_io_ipinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_54_io_ipinSE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_54_io_opinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_54_io_itrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_54_io_otrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_54_io_itrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_54_io_otrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_54_io_itrackS_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_54_io_otrackS_0; // @[CGRA.scala 273:21]
  wire  gibs_55_clock; // @[CGRA.scala 273:21]
  wire  gibs_55_reset; // @[CGRA.scala 273:21]
  wire  gibs_55_io_cfg_en; // @[CGRA.scala 273:21]
  wire [11:0] gibs_55_io_cfg_addr; // @[CGRA.scala 273:21]
  wire [31:0] gibs_55_io_cfg_data; // @[CGRA.scala 273:21]
  wire [31:0] gibs_55_io_ipinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_55_io_ipinNW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_55_io_opinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_55_io_ipinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_55_io_ipinNE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_55_io_opinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_55_io_ipinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_55_io_ipinSE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_55_io_opinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_55_io_ipinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_55_io_ipinSW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_55_io_opinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_55_io_itrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_55_io_otrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_55_io_itrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_55_io_otrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_55_io_itrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_55_io_otrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_55_io_itrackS_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_55_io_otrackS_0; // @[CGRA.scala 273:21]
  wire  gibs_56_clock; // @[CGRA.scala 273:21]
  wire  gibs_56_reset; // @[CGRA.scala 273:21]
  wire  gibs_56_io_cfg_en; // @[CGRA.scala 273:21]
  wire [11:0] gibs_56_io_cfg_addr; // @[CGRA.scala 273:21]
  wire [31:0] gibs_56_io_cfg_data; // @[CGRA.scala 273:21]
  wire [31:0] gibs_56_io_ipinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_56_io_ipinNW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_56_io_opinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_56_io_ipinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_56_io_ipinNE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_56_io_opinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_56_io_ipinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_56_io_ipinSE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_56_io_opinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_56_io_ipinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_56_io_ipinSW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_56_io_opinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_56_io_itrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_56_io_otrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_56_io_itrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_56_io_otrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_56_io_itrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_56_io_otrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_56_io_itrackS_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_56_io_otrackS_0; // @[CGRA.scala 273:21]
  wire  gibs_57_clock; // @[CGRA.scala 273:21]
  wire  gibs_57_reset; // @[CGRA.scala 273:21]
  wire  gibs_57_io_cfg_en; // @[CGRA.scala 273:21]
  wire [11:0] gibs_57_io_cfg_addr; // @[CGRA.scala 273:21]
  wire [31:0] gibs_57_io_cfg_data; // @[CGRA.scala 273:21]
  wire [31:0] gibs_57_io_ipinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_57_io_ipinNW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_57_io_opinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_57_io_ipinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_57_io_ipinNE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_57_io_opinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_57_io_ipinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_57_io_ipinSE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_57_io_opinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_57_io_ipinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_57_io_ipinSW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_57_io_opinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_57_io_itrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_57_io_otrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_57_io_itrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_57_io_otrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_57_io_itrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_57_io_otrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_57_io_itrackS_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_57_io_otrackS_0; // @[CGRA.scala 273:21]
  wire  gibs_58_clock; // @[CGRA.scala 273:21]
  wire  gibs_58_reset; // @[CGRA.scala 273:21]
  wire  gibs_58_io_cfg_en; // @[CGRA.scala 273:21]
  wire [11:0] gibs_58_io_cfg_addr; // @[CGRA.scala 273:21]
  wire [31:0] gibs_58_io_cfg_data; // @[CGRA.scala 273:21]
  wire [31:0] gibs_58_io_ipinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_58_io_ipinNW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_58_io_opinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_58_io_ipinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_58_io_ipinNE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_58_io_opinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_58_io_ipinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_58_io_ipinSE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_58_io_opinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_58_io_ipinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_58_io_ipinSW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_58_io_opinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_58_io_itrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_58_io_otrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_58_io_itrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_58_io_otrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_58_io_itrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_58_io_otrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_58_io_itrackS_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_58_io_otrackS_0; // @[CGRA.scala 273:21]
  wire  gibs_59_clock; // @[CGRA.scala 273:21]
  wire  gibs_59_reset; // @[CGRA.scala 273:21]
  wire  gibs_59_io_cfg_en; // @[CGRA.scala 273:21]
  wire [11:0] gibs_59_io_cfg_addr; // @[CGRA.scala 273:21]
  wire [31:0] gibs_59_io_cfg_data; // @[CGRA.scala 273:21]
  wire [31:0] gibs_59_io_ipinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_59_io_ipinNW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_59_io_opinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_59_io_ipinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_59_io_ipinNE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_59_io_opinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_59_io_ipinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_59_io_ipinSE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_59_io_opinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_59_io_ipinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_59_io_ipinSW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_59_io_opinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_59_io_itrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_59_io_otrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_59_io_itrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_59_io_otrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_59_io_itrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_59_io_otrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_59_io_itrackS_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_59_io_otrackS_0; // @[CGRA.scala 273:21]
  wire  gibs_60_clock; // @[CGRA.scala 273:21]
  wire  gibs_60_reset; // @[CGRA.scala 273:21]
  wire  gibs_60_io_cfg_en; // @[CGRA.scala 273:21]
  wire [11:0] gibs_60_io_cfg_addr; // @[CGRA.scala 273:21]
  wire [31:0] gibs_60_io_cfg_data; // @[CGRA.scala 273:21]
  wire [31:0] gibs_60_io_ipinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_60_io_ipinNW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_60_io_opinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_60_io_ipinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_60_io_ipinNE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_60_io_opinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_60_io_ipinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_60_io_ipinSE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_60_io_opinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_60_io_ipinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_60_io_ipinSW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_60_io_opinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_60_io_itrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_60_io_otrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_60_io_itrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_60_io_otrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_60_io_itrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_60_io_otrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_60_io_itrackS_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_60_io_otrackS_0; // @[CGRA.scala 273:21]
  wire  gibs_61_clock; // @[CGRA.scala 273:21]
  wire  gibs_61_reset; // @[CGRA.scala 273:21]
  wire  gibs_61_io_cfg_en; // @[CGRA.scala 273:21]
  wire [11:0] gibs_61_io_cfg_addr; // @[CGRA.scala 273:21]
  wire [31:0] gibs_61_io_cfg_data; // @[CGRA.scala 273:21]
  wire [31:0] gibs_61_io_ipinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_61_io_ipinNW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_61_io_opinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_61_io_ipinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_61_io_ipinNE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_61_io_opinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_61_io_ipinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_61_io_ipinSE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_61_io_opinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_61_io_ipinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_61_io_ipinSW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_61_io_opinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_61_io_itrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_61_io_otrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_61_io_itrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_61_io_otrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_61_io_itrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_61_io_otrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_61_io_itrackS_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_61_io_otrackS_0; // @[CGRA.scala 273:21]
  wire  gibs_62_clock; // @[CGRA.scala 273:21]
  wire  gibs_62_reset; // @[CGRA.scala 273:21]
  wire  gibs_62_io_cfg_en; // @[CGRA.scala 273:21]
  wire [11:0] gibs_62_io_cfg_addr; // @[CGRA.scala 273:21]
  wire [31:0] gibs_62_io_cfg_data; // @[CGRA.scala 273:21]
  wire [31:0] gibs_62_io_ipinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_62_io_ipinNW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_62_io_opinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_62_io_ipinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_62_io_ipinSW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_62_io_opinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_62_io_itrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_62_io_otrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_62_io_itrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_62_io_otrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_62_io_itrackS_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_62_io_otrackS_0; // @[CGRA.scala 273:21]
  wire  gibs_63_clock; // @[CGRA.scala 273:21]
  wire  gibs_63_reset; // @[CGRA.scala 273:21]
  wire  gibs_63_io_cfg_en; // @[CGRA.scala 273:21]
  wire [11:0] gibs_63_io_cfg_addr; // @[CGRA.scala 273:21]
  wire [31:0] gibs_63_io_cfg_data; // @[CGRA.scala 273:21]
  wire [31:0] gibs_63_io_ipinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_63_io_ipinNE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_63_io_opinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_63_io_ipinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_63_io_ipinSE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_63_io_opinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_63_io_itrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_63_io_otrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_63_io_itrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_63_io_otrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_63_io_itrackS_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_63_io_otrackS_0; // @[CGRA.scala 273:21]
  wire  gibs_64_clock; // @[CGRA.scala 273:21]
  wire  gibs_64_reset; // @[CGRA.scala 273:21]
  wire  gibs_64_io_cfg_en; // @[CGRA.scala 273:21]
  wire [11:0] gibs_64_io_cfg_addr; // @[CGRA.scala 273:21]
  wire [31:0] gibs_64_io_cfg_data; // @[CGRA.scala 273:21]
  wire [31:0] gibs_64_io_ipinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_64_io_ipinNW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_64_io_opinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_64_io_ipinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_64_io_ipinNE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_64_io_opinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_64_io_ipinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_64_io_ipinSE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_64_io_opinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_64_io_ipinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_64_io_ipinSW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_64_io_opinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_64_io_itrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_64_io_otrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_64_io_itrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_64_io_otrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_64_io_itrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_64_io_otrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_64_io_itrackS_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_64_io_otrackS_0; // @[CGRA.scala 273:21]
  wire  gibs_65_clock; // @[CGRA.scala 273:21]
  wire  gibs_65_reset; // @[CGRA.scala 273:21]
  wire  gibs_65_io_cfg_en; // @[CGRA.scala 273:21]
  wire [11:0] gibs_65_io_cfg_addr; // @[CGRA.scala 273:21]
  wire [31:0] gibs_65_io_cfg_data; // @[CGRA.scala 273:21]
  wire [31:0] gibs_65_io_ipinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_65_io_ipinNW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_65_io_opinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_65_io_ipinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_65_io_ipinNE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_65_io_opinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_65_io_ipinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_65_io_ipinSE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_65_io_opinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_65_io_ipinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_65_io_ipinSW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_65_io_opinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_65_io_itrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_65_io_otrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_65_io_itrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_65_io_otrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_65_io_itrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_65_io_otrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_65_io_itrackS_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_65_io_otrackS_0; // @[CGRA.scala 273:21]
  wire  gibs_66_clock; // @[CGRA.scala 273:21]
  wire  gibs_66_reset; // @[CGRA.scala 273:21]
  wire  gibs_66_io_cfg_en; // @[CGRA.scala 273:21]
  wire [11:0] gibs_66_io_cfg_addr; // @[CGRA.scala 273:21]
  wire [31:0] gibs_66_io_cfg_data; // @[CGRA.scala 273:21]
  wire [31:0] gibs_66_io_ipinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_66_io_ipinNW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_66_io_opinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_66_io_ipinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_66_io_ipinNE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_66_io_opinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_66_io_ipinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_66_io_ipinSE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_66_io_opinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_66_io_ipinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_66_io_ipinSW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_66_io_opinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_66_io_itrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_66_io_otrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_66_io_itrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_66_io_otrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_66_io_itrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_66_io_otrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_66_io_itrackS_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_66_io_otrackS_0; // @[CGRA.scala 273:21]
  wire  gibs_67_clock; // @[CGRA.scala 273:21]
  wire  gibs_67_reset; // @[CGRA.scala 273:21]
  wire  gibs_67_io_cfg_en; // @[CGRA.scala 273:21]
  wire [11:0] gibs_67_io_cfg_addr; // @[CGRA.scala 273:21]
  wire [31:0] gibs_67_io_cfg_data; // @[CGRA.scala 273:21]
  wire [31:0] gibs_67_io_ipinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_67_io_ipinNW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_67_io_opinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_67_io_ipinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_67_io_ipinNE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_67_io_opinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_67_io_ipinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_67_io_ipinSE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_67_io_opinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_67_io_ipinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_67_io_ipinSW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_67_io_opinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_67_io_itrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_67_io_otrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_67_io_itrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_67_io_otrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_67_io_itrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_67_io_otrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_67_io_itrackS_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_67_io_otrackS_0; // @[CGRA.scala 273:21]
  wire  gibs_68_clock; // @[CGRA.scala 273:21]
  wire  gibs_68_reset; // @[CGRA.scala 273:21]
  wire  gibs_68_io_cfg_en; // @[CGRA.scala 273:21]
  wire [11:0] gibs_68_io_cfg_addr; // @[CGRA.scala 273:21]
  wire [31:0] gibs_68_io_cfg_data; // @[CGRA.scala 273:21]
  wire [31:0] gibs_68_io_ipinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_68_io_ipinNW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_68_io_opinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_68_io_ipinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_68_io_ipinNE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_68_io_opinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_68_io_ipinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_68_io_ipinSE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_68_io_opinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_68_io_ipinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_68_io_ipinSW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_68_io_opinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_68_io_itrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_68_io_otrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_68_io_itrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_68_io_otrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_68_io_itrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_68_io_otrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_68_io_itrackS_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_68_io_otrackS_0; // @[CGRA.scala 273:21]
  wire  gibs_69_clock; // @[CGRA.scala 273:21]
  wire  gibs_69_reset; // @[CGRA.scala 273:21]
  wire  gibs_69_io_cfg_en; // @[CGRA.scala 273:21]
  wire [11:0] gibs_69_io_cfg_addr; // @[CGRA.scala 273:21]
  wire [31:0] gibs_69_io_cfg_data; // @[CGRA.scala 273:21]
  wire [31:0] gibs_69_io_ipinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_69_io_ipinNW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_69_io_opinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_69_io_ipinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_69_io_ipinNE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_69_io_opinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_69_io_ipinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_69_io_ipinSE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_69_io_opinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_69_io_ipinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_69_io_ipinSW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_69_io_opinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_69_io_itrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_69_io_otrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_69_io_itrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_69_io_otrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_69_io_itrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_69_io_otrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_69_io_itrackS_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_69_io_otrackS_0; // @[CGRA.scala 273:21]
  wire  gibs_70_clock; // @[CGRA.scala 273:21]
  wire  gibs_70_reset; // @[CGRA.scala 273:21]
  wire  gibs_70_io_cfg_en; // @[CGRA.scala 273:21]
  wire [11:0] gibs_70_io_cfg_addr; // @[CGRA.scala 273:21]
  wire [31:0] gibs_70_io_cfg_data; // @[CGRA.scala 273:21]
  wire [31:0] gibs_70_io_ipinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_70_io_ipinNW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_70_io_opinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_70_io_ipinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_70_io_ipinNE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_70_io_opinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_70_io_ipinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_70_io_ipinSE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_70_io_opinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_70_io_ipinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_70_io_ipinSW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_70_io_opinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_70_io_itrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_70_io_otrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_70_io_itrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_70_io_otrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_70_io_itrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_70_io_otrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_70_io_itrackS_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_70_io_otrackS_0; // @[CGRA.scala 273:21]
  wire  gibs_71_clock; // @[CGRA.scala 273:21]
  wire  gibs_71_reset; // @[CGRA.scala 273:21]
  wire  gibs_71_io_cfg_en; // @[CGRA.scala 273:21]
  wire [11:0] gibs_71_io_cfg_addr; // @[CGRA.scala 273:21]
  wire [31:0] gibs_71_io_cfg_data; // @[CGRA.scala 273:21]
  wire [31:0] gibs_71_io_ipinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_71_io_ipinNW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_71_io_opinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_71_io_ipinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_71_io_ipinSW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_71_io_opinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_71_io_itrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_71_io_otrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_71_io_itrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_71_io_otrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_71_io_itrackS_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_71_io_otrackS_0; // @[CGRA.scala 273:21]
  wire  gibs_72_clock; // @[CGRA.scala 273:21]
  wire  gibs_72_reset; // @[CGRA.scala 273:21]
  wire  gibs_72_io_cfg_en; // @[CGRA.scala 273:21]
  wire [11:0] gibs_72_io_cfg_addr; // @[CGRA.scala 273:21]
  wire [31:0] gibs_72_io_cfg_data; // @[CGRA.scala 273:21]
  wire [31:0] gibs_72_io_ipinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_72_io_ipinNE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_72_io_opinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_72_io_ipinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_72_io_opinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_72_io_itrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_72_io_otrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_72_io_itrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_72_io_otrackE_0; // @[CGRA.scala 273:21]
  wire  gibs_73_clock; // @[CGRA.scala 273:21]
  wire  gibs_73_reset; // @[CGRA.scala 273:21]
  wire  gibs_73_io_cfg_en; // @[CGRA.scala 273:21]
  wire [11:0] gibs_73_io_cfg_addr; // @[CGRA.scala 273:21]
  wire [31:0] gibs_73_io_cfg_data; // @[CGRA.scala 273:21]
  wire [31:0] gibs_73_io_ipinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_73_io_ipinNW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_73_io_opinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_73_io_ipinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_73_io_ipinNE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_73_io_opinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_73_io_ipinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_73_io_opinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_73_io_ipinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_73_io_opinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_73_io_itrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_73_io_otrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_73_io_itrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_73_io_otrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_73_io_itrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_73_io_otrackE_0; // @[CGRA.scala 273:21]
  wire  gibs_74_clock; // @[CGRA.scala 273:21]
  wire  gibs_74_reset; // @[CGRA.scala 273:21]
  wire  gibs_74_io_cfg_en; // @[CGRA.scala 273:21]
  wire [11:0] gibs_74_io_cfg_addr; // @[CGRA.scala 273:21]
  wire [31:0] gibs_74_io_cfg_data; // @[CGRA.scala 273:21]
  wire [31:0] gibs_74_io_ipinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_74_io_ipinNW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_74_io_opinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_74_io_ipinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_74_io_ipinNE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_74_io_opinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_74_io_ipinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_74_io_opinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_74_io_ipinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_74_io_opinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_74_io_itrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_74_io_otrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_74_io_itrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_74_io_otrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_74_io_itrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_74_io_otrackE_0; // @[CGRA.scala 273:21]
  wire  gibs_75_clock; // @[CGRA.scala 273:21]
  wire  gibs_75_reset; // @[CGRA.scala 273:21]
  wire  gibs_75_io_cfg_en; // @[CGRA.scala 273:21]
  wire [11:0] gibs_75_io_cfg_addr; // @[CGRA.scala 273:21]
  wire [31:0] gibs_75_io_cfg_data; // @[CGRA.scala 273:21]
  wire [31:0] gibs_75_io_ipinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_75_io_ipinNW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_75_io_opinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_75_io_ipinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_75_io_ipinNE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_75_io_opinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_75_io_ipinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_75_io_opinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_75_io_ipinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_75_io_opinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_75_io_itrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_75_io_otrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_75_io_itrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_75_io_otrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_75_io_itrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_75_io_otrackE_0; // @[CGRA.scala 273:21]
  wire  gibs_76_clock; // @[CGRA.scala 273:21]
  wire  gibs_76_reset; // @[CGRA.scala 273:21]
  wire  gibs_76_io_cfg_en; // @[CGRA.scala 273:21]
  wire [11:0] gibs_76_io_cfg_addr; // @[CGRA.scala 273:21]
  wire [31:0] gibs_76_io_cfg_data; // @[CGRA.scala 273:21]
  wire [31:0] gibs_76_io_ipinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_76_io_ipinNW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_76_io_opinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_76_io_ipinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_76_io_ipinNE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_76_io_opinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_76_io_ipinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_76_io_opinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_76_io_ipinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_76_io_opinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_76_io_itrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_76_io_otrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_76_io_itrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_76_io_otrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_76_io_itrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_76_io_otrackE_0; // @[CGRA.scala 273:21]
  wire  gibs_77_clock; // @[CGRA.scala 273:21]
  wire  gibs_77_reset; // @[CGRA.scala 273:21]
  wire  gibs_77_io_cfg_en; // @[CGRA.scala 273:21]
  wire [11:0] gibs_77_io_cfg_addr; // @[CGRA.scala 273:21]
  wire [31:0] gibs_77_io_cfg_data; // @[CGRA.scala 273:21]
  wire [31:0] gibs_77_io_ipinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_77_io_ipinNW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_77_io_opinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_77_io_ipinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_77_io_ipinNE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_77_io_opinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_77_io_ipinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_77_io_opinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_77_io_ipinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_77_io_opinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_77_io_itrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_77_io_otrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_77_io_itrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_77_io_otrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_77_io_itrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_77_io_otrackE_0; // @[CGRA.scala 273:21]
  wire  gibs_78_clock; // @[CGRA.scala 273:21]
  wire  gibs_78_reset; // @[CGRA.scala 273:21]
  wire  gibs_78_io_cfg_en; // @[CGRA.scala 273:21]
  wire [11:0] gibs_78_io_cfg_addr; // @[CGRA.scala 273:21]
  wire [31:0] gibs_78_io_cfg_data; // @[CGRA.scala 273:21]
  wire [31:0] gibs_78_io_ipinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_78_io_ipinNW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_78_io_opinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_78_io_ipinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_78_io_ipinNE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_78_io_opinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_78_io_ipinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_78_io_opinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_78_io_ipinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_78_io_opinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_78_io_itrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_78_io_otrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_78_io_itrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_78_io_otrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_78_io_itrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_78_io_otrackE_0; // @[CGRA.scala 273:21]
  wire  gibs_79_clock; // @[CGRA.scala 273:21]
  wire  gibs_79_reset; // @[CGRA.scala 273:21]
  wire  gibs_79_io_cfg_en; // @[CGRA.scala 273:21]
  wire [11:0] gibs_79_io_cfg_addr; // @[CGRA.scala 273:21]
  wire [31:0] gibs_79_io_cfg_data; // @[CGRA.scala 273:21]
  wire [31:0] gibs_79_io_ipinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_79_io_ipinNW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_79_io_opinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_79_io_ipinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_79_io_ipinNE_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_79_io_opinNE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_79_io_ipinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_79_io_opinSE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_79_io_ipinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_79_io_opinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_79_io_itrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_79_io_otrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_79_io_itrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_79_io_otrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_79_io_itrackE_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_79_io_otrackE_0; // @[CGRA.scala 273:21]
  wire  gibs_80_clock; // @[CGRA.scala 273:21]
  wire  gibs_80_reset; // @[CGRA.scala 273:21]
  wire  gibs_80_io_cfg_en; // @[CGRA.scala 273:21]
  wire [11:0] gibs_80_io_cfg_addr; // @[CGRA.scala 273:21]
  wire [31:0] gibs_80_io_cfg_data; // @[CGRA.scala 273:21]
  wire [31:0] gibs_80_io_ipinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_80_io_ipinNW_1; // @[CGRA.scala 273:21]
  wire [31:0] gibs_80_io_opinNW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_80_io_ipinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_80_io_opinSW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_80_io_itrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_80_io_otrackW_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_80_io_itrackN_0; // @[CGRA.scala 273:21]
  wire [31:0] gibs_80_io_otrackN_0; // @[CGRA.scala 273:21]
  reg [44:0] cfgRegs_0; // @[CGRA.scala 487:24]
  reg [44:0] cfgRegs_1; // @[CGRA.scala 487:24]
  reg [44:0] cfgRegs_2; // @[CGRA.scala 487:24]
  reg [44:0] cfgRegs_3; // @[CGRA.scala 487:24]
  reg [44:0] cfgRegs_4; // @[CGRA.scala 487:24]
  reg [44:0] cfgRegs_5; // @[CGRA.scala 487:24]
  reg [44:0] cfgRegs_6; // @[CGRA.scala 487:24]
  reg [44:0] cfgRegs_7; // @[CGRA.scala 487:24]
  reg [44:0] cfgRegs_8; // @[CGRA.scala 487:24]
  reg [44:0] cfgRegs_9; // @[CGRA.scala 487:24]
  reg [44:0] cfgRegs_10; // @[CGRA.scala 487:24]
  reg [44:0] cfgRegs_11; // @[CGRA.scala 487:24]
  reg [44:0] cfgRegs_12; // @[CGRA.scala 487:24]
  reg [44:0] cfgRegs_13; // @[CGRA.scala 487:24]
  reg [44:0] cfgRegs_14; // @[CGRA.scala 487:24]
  reg [44:0] cfgRegs_15; // @[CGRA.scala 487:24]
  reg [44:0] cfgRegs_16; // @[CGRA.scala 487:24]
  reg [44:0] cfgRegs_17; // @[CGRA.scala 487:24]
  reg [44:0] cfgRegs_18; // @[CGRA.scala 487:24]
  reg [44:0] cfgRegs_19; // @[CGRA.scala 487:24]
  wire [44:0] _T_2 = {io_cfg_en,io_cfg_addr,io_cfg_data}; // @[Cat.scala 29:58]
  IOB ibs_0 ( // @[CGRA.scala 149:20]
    .io_in_0(ibs_0_io_in_0),
    .io_out_0(ibs_0_io_out_0)
  );
  IOB ibs_1 ( // @[CGRA.scala 149:20]
    .io_in_0(ibs_1_io_in_0),
    .io_out_0(ibs_1_io_out_0)
  );
  IOB ibs_2 ( // @[CGRA.scala 149:20]
    .io_in_0(ibs_2_io_in_0),
    .io_out_0(ibs_2_io_out_0)
  );
  IOB ibs_3 ( // @[CGRA.scala 149:20]
    .io_in_0(ibs_3_io_in_0),
    .io_out_0(ibs_3_io_out_0)
  );
  IOB ibs_4 ( // @[CGRA.scala 149:20]
    .io_in_0(ibs_4_io_in_0),
    .io_out_0(ibs_4_io_out_0)
  );
  IOB ibs_5 ( // @[CGRA.scala 149:20]
    .io_in_0(ibs_5_io_in_0),
    .io_out_0(ibs_5_io_out_0)
  );
  IOB ibs_6 ( // @[CGRA.scala 149:20]
    .io_in_0(ibs_6_io_in_0),
    .io_out_0(ibs_6_io_out_0)
  );
  IOB ibs_7 ( // @[CGRA.scala 149:20]
    .io_in_0(ibs_7_io_in_0),
    .io_out_0(ibs_7_io_out_0)
  );
  IOB ibs_8 ( // @[CGRA.scala 149:20]
    .io_in_0(ibs_8_io_in_0),
    .io_out_0(ibs_8_io_out_0)
  );
  IOB ibs_9 ( // @[CGRA.scala 149:20]
    .io_in_0(ibs_9_io_in_0),
    .io_out_0(ibs_9_io_out_0)
  );
  IOB ibs_10 ( // @[CGRA.scala 149:20]
    .io_in_0(ibs_10_io_in_0),
    .io_out_0(ibs_10_io_out_0)
  );
  IOB ibs_11 ( // @[CGRA.scala 149:20]
    .io_in_0(ibs_11_io_in_0),
    .io_out_0(ibs_11_io_out_0)
  );
  IOB ibs_12 ( // @[CGRA.scala 149:20]
    .io_in_0(ibs_12_io_in_0),
    .io_out_0(ibs_12_io_out_0)
  );
  IOB ibs_13 ( // @[CGRA.scala 149:20]
    .io_in_0(ibs_13_io_in_0),
    .io_out_0(ibs_13_io_out_0)
  );
  IOB ibs_14 ( // @[CGRA.scala 149:20]
    .io_in_0(ibs_14_io_in_0),
    .io_out_0(ibs_14_io_out_0)
  );
  IOB ibs_15 ( // @[CGRA.scala 149:20]
    .io_in_0(ibs_15_io_in_0),
    .io_out_0(ibs_15_io_out_0)
  );
  IOB_16 obs_0 ( // @[CGRA.scala 176:20]
    .clock(obs_0_clock),
    .reset(obs_0_reset),
    .io_cfg_en(obs_0_io_cfg_en),
    .io_cfg_addr(obs_0_io_cfg_addr),
    .io_cfg_data(obs_0_io_cfg_data),
    .io_in_0(obs_0_io_in_0),
    .io_in_1(obs_0_io_in_1),
    .io_out_0(obs_0_io_out_0)
  );
  IOB_17 obs_1 ( // @[CGRA.scala 176:20]
    .clock(obs_1_clock),
    .reset(obs_1_reset),
    .io_cfg_en(obs_1_io_cfg_en),
    .io_cfg_addr(obs_1_io_cfg_addr),
    .io_cfg_data(obs_1_io_cfg_data),
    .io_in_0(obs_1_io_in_0),
    .io_in_1(obs_1_io_in_1),
    .io_out_0(obs_1_io_out_0)
  );
  IOB_18 obs_2 ( // @[CGRA.scala 176:20]
    .clock(obs_2_clock),
    .reset(obs_2_reset),
    .io_cfg_en(obs_2_io_cfg_en),
    .io_cfg_addr(obs_2_io_cfg_addr),
    .io_cfg_data(obs_2_io_cfg_data),
    .io_in_0(obs_2_io_in_0),
    .io_in_1(obs_2_io_in_1),
    .io_out_0(obs_2_io_out_0)
  );
  IOB_19 obs_3 ( // @[CGRA.scala 176:20]
    .clock(obs_3_clock),
    .reset(obs_3_reset),
    .io_cfg_en(obs_3_io_cfg_en),
    .io_cfg_addr(obs_3_io_cfg_addr),
    .io_cfg_data(obs_3_io_cfg_data),
    .io_in_0(obs_3_io_in_0),
    .io_in_1(obs_3_io_in_1),
    .io_out_0(obs_3_io_out_0)
  );
  IOB_20 obs_4 ( // @[CGRA.scala 176:20]
    .clock(obs_4_clock),
    .reset(obs_4_reset),
    .io_cfg_en(obs_4_io_cfg_en),
    .io_cfg_addr(obs_4_io_cfg_addr),
    .io_cfg_data(obs_4_io_cfg_data),
    .io_in_0(obs_4_io_in_0),
    .io_in_1(obs_4_io_in_1),
    .io_out_0(obs_4_io_out_0)
  );
  IOB_21 obs_5 ( // @[CGRA.scala 176:20]
    .clock(obs_5_clock),
    .reset(obs_5_reset),
    .io_cfg_en(obs_5_io_cfg_en),
    .io_cfg_addr(obs_5_io_cfg_addr),
    .io_cfg_data(obs_5_io_cfg_data),
    .io_in_0(obs_5_io_in_0),
    .io_in_1(obs_5_io_in_1),
    .io_out_0(obs_5_io_out_0)
  );
  IOB_22 obs_6 ( // @[CGRA.scala 176:20]
    .clock(obs_6_clock),
    .reset(obs_6_reset),
    .io_cfg_en(obs_6_io_cfg_en),
    .io_cfg_addr(obs_6_io_cfg_addr),
    .io_cfg_data(obs_6_io_cfg_data),
    .io_in_0(obs_6_io_in_0),
    .io_in_1(obs_6_io_in_1),
    .io_out_0(obs_6_io_out_0)
  );
  IOB_23 obs_7 ( // @[CGRA.scala 176:20]
    .clock(obs_7_clock),
    .reset(obs_7_reset),
    .io_cfg_en(obs_7_io_cfg_en),
    .io_cfg_addr(obs_7_io_cfg_addr),
    .io_cfg_data(obs_7_io_cfg_data),
    .io_in_0(obs_7_io_in_0),
    .io_in_1(obs_7_io_in_1),
    .io_out_0(obs_7_io_out_0)
  );
  IOB_24 obs_8 ( // @[CGRA.scala 176:20]
    .clock(obs_8_clock),
    .reset(obs_8_reset),
    .io_cfg_en(obs_8_io_cfg_en),
    .io_cfg_addr(obs_8_io_cfg_addr),
    .io_cfg_data(obs_8_io_cfg_data),
    .io_in_0(obs_8_io_in_0),
    .io_in_1(obs_8_io_in_1),
    .io_out_0(obs_8_io_out_0)
  );
  IOB_25 obs_9 ( // @[CGRA.scala 176:20]
    .clock(obs_9_clock),
    .reset(obs_9_reset),
    .io_cfg_en(obs_9_io_cfg_en),
    .io_cfg_addr(obs_9_io_cfg_addr),
    .io_cfg_data(obs_9_io_cfg_data),
    .io_in_0(obs_9_io_in_0),
    .io_in_1(obs_9_io_in_1),
    .io_out_0(obs_9_io_out_0)
  );
  IOB_26 obs_10 ( // @[CGRA.scala 176:20]
    .clock(obs_10_clock),
    .reset(obs_10_reset),
    .io_cfg_en(obs_10_io_cfg_en),
    .io_cfg_addr(obs_10_io_cfg_addr),
    .io_cfg_data(obs_10_io_cfg_data),
    .io_in_0(obs_10_io_in_0),
    .io_in_1(obs_10_io_in_1),
    .io_out_0(obs_10_io_out_0)
  );
  IOB_27 obs_11 ( // @[CGRA.scala 176:20]
    .clock(obs_11_clock),
    .reset(obs_11_reset),
    .io_cfg_en(obs_11_io_cfg_en),
    .io_cfg_addr(obs_11_io_cfg_addr),
    .io_cfg_data(obs_11_io_cfg_data),
    .io_in_0(obs_11_io_in_0),
    .io_in_1(obs_11_io_in_1),
    .io_out_0(obs_11_io_out_0)
  );
  IOB_28 obs_12 ( // @[CGRA.scala 176:20]
    .clock(obs_12_clock),
    .reset(obs_12_reset),
    .io_cfg_en(obs_12_io_cfg_en),
    .io_cfg_addr(obs_12_io_cfg_addr),
    .io_cfg_data(obs_12_io_cfg_data),
    .io_in_0(obs_12_io_in_0),
    .io_in_1(obs_12_io_in_1),
    .io_out_0(obs_12_io_out_0)
  );
  IOB_29 obs_13 ( // @[CGRA.scala 176:20]
    .clock(obs_13_clock),
    .reset(obs_13_reset),
    .io_cfg_en(obs_13_io_cfg_en),
    .io_cfg_addr(obs_13_io_cfg_addr),
    .io_cfg_data(obs_13_io_cfg_data),
    .io_in_0(obs_13_io_in_0),
    .io_in_1(obs_13_io_in_1),
    .io_out_0(obs_13_io_out_0)
  );
  IOB_30 obs_14 ( // @[CGRA.scala 176:20]
    .clock(obs_14_clock),
    .reset(obs_14_reset),
    .io_cfg_en(obs_14_io_cfg_en),
    .io_cfg_addr(obs_14_io_cfg_addr),
    .io_cfg_data(obs_14_io_cfg_data),
    .io_in_0(obs_14_io_in_0),
    .io_in_1(obs_14_io_in_1),
    .io_out_0(obs_14_io_out_0)
  );
  IOB_31 obs_15 ( // @[CGRA.scala 176:20]
    .clock(obs_15_clock),
    .reset(obs_15_reset),
    .io_cfg_en(obs_15_io_cfg_en),
    .io_cfg_addr(obs_15_io_cfg_addr),
    .io_cfg_data(obs_15_io_cfg_data),
    .io_in_0(obs_15_io_in_0),
    .io_in_1(obs_15_io_in_1),
    .io_out_0(obs_15_io_out_0)
  );
  GPE pes_0 ( // @[CGRA.scala 200:20]
    .clock(pes_0_clock),
    .reset(pes_0_reset),
    .io_cfg_en(pes_0_io_cfg_en),
    .io_cfg_addr(pes_0_io_cfg_addr),
    .io_cfg_data(pes_0_io_cfg_data),
    .io_en(pes_0_io_en),
    .io_in_0(pes_0_io_in_0),
    .io_in_1(pes_0_io_in_1),
    .io_in_2(pes_0_io_in_2),
    .io_in_3(pes_0_io_in_3),
    .io_in_4(pes_0_io_in_4),
    .io_in_5(pes_0_io_in_5),
    .io_in_6(pes_0_io_in_6),
    .io_in_7(pes_0_io_in_7),
    .io_out_0(pes_0_io_out_0)
  );
  GPE_1 pes_1 ( // @[CGRA.scala 200:20]
    .clock(pes_1_clock),
    .reset(pes_1_reset),
    .io_cfg_en(pes_1_io_cfg_en),
    .io_cfg_addr(pes_1_io_cfg_addr),
    .io_cfg_data(pes_1_io_cfg_data),
    .io_en(pes_1_io_en),
    .io_in_0(pes_1_io_in_0),
    .io_in_1(pes_1_io_in_1),
    .io_in_2(pes_1_io_in_2),
    .io_in_3(pes_1_io_in_3),
    .io_in_4(pes_1_io_in_4),
    .io_in_5(pes_1_io_in_5),
    .io_in_6(pes_1_io_in_6),
    .io_in_7(pes_1_io_in_7),
    .io_out_0(pes_1_io_out_0)
  );
  GPE_2 pes_2 ( // @[CGRA.scala 200:20]
    .clock(pes_2_clock),
    .reset(pes_2_reset),
    .io_cfg_en(pes_2_io_cfg_en),
    .io_cfg_addr(pes_2_io_cfg_addr),
    .io_cfg_data(pes_2_io_cfg_data),
    .io_en(pes_2_io_en),
    .io_in_0(pes_2_io_in_0),
    .io_in_1(pes_2_io_in_1),
    .io_in_2(pes_2_io_in_2),
    .io_in_3(pes_2_io_in_3),
    .io_in_4(pes_2_io_in_4),
    .io_in_5(pes_2_io_in_5),
    .io_in_6(pes_2_io_in_6),
    .io_in_7(pes_2_io_in_7),
    .io_out_0(pes_2_io_out_0)
  );
  GPE_3 pes_3 ( // @[CGRA.scala 200:20]
    .clock(pes_3_clock),
    .reset(pes_3_reset),
    .io_cfg_en(pes_3_io_cfg_en),
    .io_cfg_addr(pes_3_io_cfg_addr),
    .io_cfg_data(pes_3_io_cfg_data),
    .io_en(pes_3_io_en),
    .io_in_0(pes_3_io_in_0),
    .io_in_1(pes_3_io_in_1),
    .io_in_2(pes_3_io_in_2),
    .io_in_3(pes_3_io_in_3),
    .io_in_4(pes_3_io_in_4),
    .io_in_5(pes_3_io_in_5),
    .io_in_6(pes_3_io_in_6),
    .io_in_7(pes_3_io_in_7),
    .io_out_0(pes_3_io_out_0)
  );
  GPE_4 pes_4 ( // @[CGRA.scala 200:20]
    .clock(pes_4_clock),
    .reset(pes_4_reset),
    .io_cfg_en(pes_4_io_cfg_en),
    .io_cfg_addr(pes_4_io_cfg_addr),
    .io_cfg_data(pes_4_io_cfg_data),
    .io_en(pes_4_io_en),
    .io_in_0(pes_4_io_in_0),
    .io_in_1(pes_4_io_in_1),
    .io_in_2(pes_4_io_in_2),
    .io_in_3(pes_4_io_in_3),
    .io_in_4(pes_4_io_in_4),
    .io_in_5(pes_4_io_in_5),
    .io_in_6(pes_4_io_in_6),
    .io_in_7(pes_4_io_in_7),
    .io_out_0(pes_4_io_out_0)
  );
  GPE_5 pes_5 ( // @[CGRA.scala 200:20]
    .clock(pes_5_clock),
    .reset(pes_5_reset),
    .io_cfg_en(pes_5_io_cfg_en),
    .io_cfg_addr(pes_5_io_cfg_addr),
    .io_cfg_data(pes_5_io_cfg_data),
    .io_en(pes_5_io_en),
    .io_in_0(pes_5_io_in_0),
    .io_in_1(pes_5_io_in_1),
    .io_in_2(pes_5_io_in_2),
    .io_in_3(pes_5_io_in_3),
    .io_in_4(pes_5_io_in_4),
    .io_in_5(pes_5_io_in_5),
    .io_in_6(pes_5_io_in_6),
    .io_in_7(pes_5_io_in_7),
    .io_out_0(pes_5_io_out_0)
  );
  GPE_6 pes_6 ( // @[CGRA.scala 200:20]
    .clock(pes_6_clock),
    .reset(pes_6_reset),
    .io_cfg_en(pes_6_io_cfg_en),
    .io_cfg_addr(pes_6_io_cfg_addr),
    .io_cfg_data(pes_6_io_cfg_data),
    .io_en(pes_6_io_en),
    .io_in_0(pes_6_io_in_0),
    .io_in_1(pes_6_io_in_1),
    .io_in_2(pes_6_io_in_2),
    .io_in_3(pes_6_io_in_3),
    .io_in_4(pes_6_io_in_4),
    .io_in_5(pes_6_io_in_5),
    .io_in_6(pes_6_io_in_6),
    .io_in_7(pes_6_io_in_7),
    .io_out_0(pes_6_io_out_0)
  );
  GPE_7 pes_7 ( // @[CGRA.scala 200:20]
    .clock(pes_7_clock),
    .reset(pes_7_reset),
    .io_cfg_en(pes_7_io_cfg_en),
    .io_cfg_addr(pes_7_io_cfg_addr),
    .io_cfg_data(pes_7_io_cfg_data),
    .io_en(pes_7_io_en),
    .io_in_0(pes_7_io_in_0),
    .io_in_1(pes_7_io_in_1),
    .io_in_2(pes_7_io_in_2),
    .io_in_3(pes_7_io_in_3),
    .io_in_4(pes_7_io_in_4),
    .io_in_5(pes_7_io_in_5),
    .io_in_6(pes_7_io_in_6),
    .io_in_7(pes_7_io_in_7),
    .io_out_0(pes_7_io_out_0)
  );
  GPE_8 pes_8 ( // @[CGRA.scala 200:20]
    .clock(pes_8_clock),
    .reset(pes_8_reset),
    .io_cfg_en(pes_8_io_cfg_en),
    .io_cfg_addr(pes_8_io_cfg_addr),
    .io_cfg_data(pes_8_io_cfg_data),
    .io_en(pes_8_io_en),
    .io_in_0(pes_8_io_in_0),
    .io_in_1(pes_8_io_in_1),
    .io_in_2(pes_8_io_in_2),
    .io_in_3(pes_8_io_in_3),
    .io_in_4(pes_8_io_in_4),
    .io_in_5(pes_8_io_in_5),
    .io_in_6(pes_8_io_in_6),
    .io_in_7(pes_8_io_in_7),
    .io_out_0(pes_8_io_out_0)
  );
  GPE_9 pes_9 ( // @[CGRA.scala 200:20]
    .clock(pes_9_clock),
    .reset(pes_9_reset),
    .io_cfg_en(pes_9_io_cfg_en),
    .io_cfg_addr(pes_9_io_cfg_addr),
    .io_cfg_data(pes_9_io_cfg_data),
    .io_en(pes_9_io_en),
    .io_in_0(pes_9_io_in_0),
    .io_in_1(pes_9_io_in_1),
    .io_in_2(pes_9_io_in_2),
    .io_in_3(pes_9_io_in_3),
    .io_in_4(pes_9_io_in_4),
    .io_in_5(pes_9_io_in_5),
    .io_in_6(pes_9_io_in_6),
    .io_in_7(pes_9_io_in_7),
    .io_out_0(pes_9_io_out_0)
  );
  GPE_10 pes_10 ( // @[CGRA.scala 200:20]
    .clock(pes_10_clock),
    .reset(pes_10_reset),
    .io_cfg_en(pes_10_io_cfg_en),
    .io_cfg_addr(pes_10_io_cfg_addr),
    .io_cfg_data(pes_10_io_cfg_data),
    .io_en(pes_10_io_en),
    .io_in_0(pes_10_io_in_0),
    .io_in_1(pes_10_io_in_1),
    .io_in_2(pes_10_io_in_2),
    .io_in_3(pes_10_io_in_3),
    .io_in_4(pes_10_io_in_4),
    .io_in_5(pes_10_io_in_5),
    .io_in_6(pes_10_io_in_6),
    .io_in_7(pes_10_io_in_7),
    .io_out_0(pes_10_io_out_0)
  );
  GPE_11 pes_11 ( // @[CGRA.scala 200:20]
    .clock(pes_11_clock),
    .reset(pes_11_reset),
    .io_cfg_en(pes_11_io_cfg_en),
    .io_cfg_addr(pes_11_io_cfg_addr),
    .io_cfg_data(pes_11_io_cfg_data),
    .io_en(pes_11_io_en),
    .io_in_0(pes_11_io_in_0),
    .io_in_1(pes_11_io_in_1),
    .io_in_2(pes_11_io_in_2),
    .io_in_3(pes_11_io_in_3),
    .io_in_4(pes_11_io_in_4),
    .io_in_5(pes_11_io_in_5),
    .io_in_6(pes_11_io_in_6),
    .io_in_7(pes_11_io_in_7),
    .io_out_0(pes_11_io_out_0)
  );
  GPE_12 pes_12 ( // @[CGRA.scala 200:20]
    .clock(pes_12_clock),
    .reset(pes_12_reset),
    .io_cfg_en(pes_12_io_cfg_en),
    .io_cfg_addr(pes_12_io_cfg_addr),
    .io_cfg_data(pes_12_io_cfg_data),
    .io_en(pes_12_io_en),
    .io_in_0(pes_12_io_in_0),
    .io_in_1(pes_12_io_in_1),
    .io_in_2(pes_12_io_in_2),
    .io_in_3(pes_12_io_in_3),
    .io_in_4(pes_12_io_in_4),
    .io_in_5(pes_12_io_in_5),
    .io_in_6(pes_12_io_in_6),
    .io_in_7(pes_12_io_in_7),
    .io_out_0(pes_12_io_out_0)
  );
  GPE_13 pes_13 ( // @[CGRA.scala 200:20]
    .clock(pes_13_clock),
    .reset(pes_13_reset),
    .io_cfg_en(pes_13_io_cfg_en),
    .io_cfg_addr(pes_13_io_cfg_addr),
    .io_cfg_data(pes_13_io_cfg_data),
    .io_en(pes_13_io_en),
    .io_in_0(pes_13_io_in_0),
    .io_in_1(pes_13_io_in_1),
    .io_in_2(pes_13_io_in_2),
    .io_in_3(pes_13_io_in_3),
    .io_in_4(pes_13_io_in_4),
    .io_in_5(pes_13_io_in_5),
    .io_in_6(pes_13_io_in_6),
    .io_in_7(pes_13_io_in_7),
    .io_out_0(pes_13_io_out_0)
  );
  GPE_14 pes_14 ( // @[CGRA.scala 200:20]
    .clock(pes_14_clock),
    .reset(pes_14_reset),
    .io_cfg_en(pes_14_io_cfg_en),
    .io_cfg_addr(pes_14_io_cfg_addr),
    .io_cfg_data(pes_14_io_cfg_data),
    .io_en(pes_14_io_en),
    .io_in_0(pes_14_io_in_0),
    .io_in_1(pes_14_io_in_1),
    .io_in_2(pes_14_io_in_2),
    .io_in_3(pes_14_io_in_3),
    .io_in_4(pes_14_io_in_4),
    .io_in_5(pes_14_io_in_5),
    .io_in_6(pes_14_io_in_6),
    .io_in_7(pes_14_io_in_7),
    .io_out_0(pes_14_io_out_0)
  );
  GPE_15 pes_15 ( // @[CGRA.scala 200:20]
    .clock(pes_15_clock),
    .reset(pes_15_reset),
    .io_cfg_en(pes_15_io_cfg_en),
    .io_cfg_addr(pes_15_io_cfg_addr),
    .io_cfg_data(pes_15_io_cfg_data),
    .io_en(pes_15_io_en),
    .io_in_0(pes_15_io_in_0),
    .io_in_1(pes_15_io_in_1),
    .io_in_2(pes_15_io_in_2),
    .io_in_3(pes_15_io_in_3),
    .io_in_4(pes_15_io_in_4),
    .io_in_5(pes_15_io_in_5),
    .io_in_6(pes_15_io_in_6),
    .io_in_7(pes_15_io_in_7),
    .io_out_0(pes_15_io_out_0)
  );
  GPE_16 pes_16 ( // @[CGRA.scala 200:20]
    .clock(pes_16_clock),
    .reset(pes_16_reset),
    .io_cfg_en(pes_16_io_cfg_en),
    .io_cfg_addr(pes_16_io_cfg_addr),
    .io_cfg_data(pes_16_io_cfg_data),
    .io_en(pes_16_io_en),
    .io_in_0(pes_16_io_in_0),
    .io_in_1(pes_16_io_in_1),
    .io_in_2(pes_16_io_in_2),
    .io_in_3(pes_16_io_in_3),
    .io_in_4(pes_16_io_in_4),
    .io_in_5(pes_16_io_in_5),
    .io_in_6(pes_16_io_in_6),
    .io_in_7(pes_16_io_in_7),
    .io_out_0(pes_16_io_out_0)
  );
  GPE_17 pes_17 ( // @[CGRA.scala 200:20]
    .clock(pes_17_clock),
    .reset(pes_17_reset),
    .io_cfg_en(pes_17_io_cfg_en),
    .io_cfg_addr(pes_17_io_cfg_addr),
    .io_cfg_data(pes_17_io_cfg_data),
    .io_en(pes_17_io_en),
    .io_in_0(pes_17_io_in_0),
    .io_in_1(pes_17_io_in_1),
    .io_in_2(pes_17_io_in_2),
    .io_in_3(pes_17_io_in_3),
    .io_in_4(pes_17_io_in_4),
    .io_in_5(pes_17_io_in_5),
    .io_in_6(pes_17_io_in_6),
    .io_in_7(pes_17_io_in_7),
    .io_out_0(pes_17_io_out_0)
  );
  GPE_18 pes_18 ( // @[CGRA.scala 200:20]
    .clock(pes_18_clock),
    .reset(pes_18_reset),
    .io_cfg_en(pes_18_io_cfg_en),
    .io_cfg_addr(pes_18_io_cfg_addr),
    .io_cfg_data(pes_18_io_cfg_data),
    .io_en(pes_18_io_en),
    .io_in_0(pes_18_io_in_0),
    .io_in_1(pes_18_io_in_1),
    .io_in_2(pes_18_io_in_2),
    .io_in_3(pes_18_io_in_3),
    .io_in_4(pes_18_io_in_4),
    .io_in_5(pes_18_io_in_5),
    .io_in_6(pes_18_io_in_6),
    .io_in_7(pes_18_io_in_7),
    .io_out_0(pes_18_io_out_0)
  );
  GPE_19 pes_19 ( // @[CGRA.scala 200:20]
    .clock(pes_19_clock),
    .reset(pes_19_reset),
    .io_cfg_en(pes_19_io_cfg_en),
    .io_cfg_addr(pes_19_io_cfg_addr),
    .io_cfg_data(pes_19_io_cfg_data),
    .io_en(pes_19_io_en),
    .io_in_0(pes_19_io_in_0),
    .io_in_1(pes_19_io_in_1),
    .io_in_2(pes_19_io_in_2),
    .io_in_3(pes_19_io_in_3),
    .io_in_4(pes_19_io_in_4),
    .io_in_5(pes_19_io_in_5),
    .io_in_6(pes_19_io_in_6),
    .io_in_7(pes_19_io_in_7),
    .io_out_0(pes_19_io_out_0)
  );
  GPE_20 pes_20 ( // @[CGRA.scala 200:20]
    .clock(pes_20_clock),
    .reset(pes_20_reset),
    .io_cfg_en(pes_20_io_cfg_en),
    .io_cfg_addr(pes_20_io_cfg_addr),
    .io_cfg_data(pes_20_io_cfg_data),
    .io_en(pes_20_io_en),
    .io_in_0(pes_20_io_in_0),
    .io_in_1(pes_20_io_in_1),
    .io_in_2(pes_20_io_in_2),
    .io_in_3(pes_20_io_in_3),
    .io_in_4(pes_20_io_in_4),
    .io_in_5(pes_20_io_in_5),
    .io_in_6(pes_20_io_in_6),
    .io_in_7(pes_20_io_in_7),
    .io_out_0(pes_20_io_out_0)
  );
  GPE_21 pes_21 ( // @[CGRA.scala 200:20]
    .clock(pes_21_clock),
    .reset(pes_21_reset),
    .io_cfg_en(pes_21_io_cfg_en),
    .io_cfg_addr(pes_21_io_cfg_addr),
    .io_cfg_data(pes_21_io_cfg_data),
    .io_en(pes_21_io_en),
    .io_in_0(pes_21_io_in_0),
    .io_in_1(pes_21_io_in_1),
    .io_in_2(pes_21_io_in_2),
    .io_in_3(pes_21_io_in_3),
    .io_in_4(pes_21_io_in_4),
    .io_in_5(pes_21_io_in_5),
    .io_in_6(pes_21_io_in_6),
    .io_in_7(pes_21_io_in_7),
    .io_out_0(pes_21_io_out_0)
  );
  GPE_22 pes_22 ( // @[CGRA.scala 200:20]
    .clock(pes_22_clock),
    .reset(pes_22_reset),
    .io_cfg_en(pes_22_io_cfg_en),
    .io_cfg_addr(pes_22_io_cfg_addr),
    .io_cfg_data(pes_22_io_cfg_data),
    .io_en(pes_22_io_en),
    .io_in_0(pes_22_io_in_0),
    .io_in_1(pes_22_io_in_1),
    .io_in_2(pes_22_io_in_2),
    .io_in_3(pes_22_io_in_3),
    .io_in_4(pes_22_io_in_4),
    .io_in_5(pes_22_io_in_5),
    .io_in_6(pes_22_io_in_6),
    .io_in_7(pes_22_io_in_7),
    .io_out_0(pes_22_io_out_0)
  );
  GPE_23 pes_23 ( // @[CGRA.scala 200:20]
    .clock(pes_23_clock),
    .reset(pes_23_reset),
    .io_cfg_en(pes_23_io_cfg_en),
    .io_cfg_addr(pes_23_io_cfg_addr),
    .io_cfg_data(pes_23_io_cfg_data),
    .io_en(pes_23_io_en),
    .io_in_0(pes_23_io_in_0),
    .io_in_1(pes_23_io_in_1),
    .io_in_2(pes_23_io_in_2),
    .io_in_3(pes_23_io_in_3),
    .io_in_4(pes_23_io_in_4),
    .io_in_5(pes_23_io_in_5),
    .io_in_6(pes_23_io_in_6),
    .io_in_7(pes_23_io_in_7),
    .io_out_0(pes_23_io_out_0)
  );
  GPE_24 pes_24 ( // @[CGRA.scala 200:20]
    .clock(pes_24_clock),
    .reset(pes_24_reset),
    .io_cfg_en(pes_24_io_cfg_en),
    .io_cfg_addr(pes_24_io_cfg_addr),
    .io_cfg_data(pes_24_io_cfg_data),
    .io_en(pes_24_io_en),
    .io_in_0(pes_24_io_in_0),
    .io_in_1(pes_24_io_in_1),
    .io_in_2(pes_24_io_in_2),
    .io_in_3(pes_24_io_in_3),
    .io_in_4(pes_24_io_in_4),
    .io_in_5(pes_24_io_in_5),
    .io_in_6(pes_24_io_in_6),
    .io_in_7(pes_24_io_in_7),
    .io_out_0(pes_24_io_out_0)
  );
  GPE_25 pes_25 ( // @[CGRA.scala 200:20]
    .clock(pes_25_clock),
    .reset(pes_25_reset),
    .io_cfg_en(pes_25_io_cfg_en),
    .io_cfg_addr(pes_25_io_cfg_addr),
    .io_cfg_data(pes_25_io_cfg_data),
    .io_en(pes_25_io_en),
    .io_in_0(pes_25_io_in_0),
    .io_in_1(pes_25_io_in_1),
    .io_in_2(pes_25_io_in_2),
    .io_in_3(pes_25_io_in_3),
    .io_in_4(pes_25_io_in_4),
    .io_in_5(pes_25_io_in_5),
    .io_in_6(pes_25_io_in_6),
    .io_in_7(pes_25_io_in_7),
    .io_out_0(pes_25_io_out_0)
  );
  GPE_26 pes_26 ( // @[CGRA.scala 200:20]
    .clock(pes_26_clock),
    .reset(pes_26_reset),
    .io_cfg_en(pes_26_io_cfg_en),
    .io_cfg_addr(pes_26_io_cfg_addr),
    .io_cfg_data(pes_26_io_cfg_data),
    .io_en(pes_26_io_en),
    .io_in_0(pes_26_io_in_0),
    .io_in_1(pes_26_io_in_1),
    .io_in_2(pes_26_io_in_2),
    .io_in_3(pes_26_io_in_3),
    .io_in_4(pes_26_io_in_4),
    .io_in_5(pes_26_io_in_5),
    .io_in_6(pes_26_io_in_6),
    .io_in_7(pes_26_io_in_7),
    .io_out_0(pes_26_io_out_0)
  );
  GPE_27 pes_27 ( // @[CGRA.scala 200:20]
    .clock(pes_27_clock),
    .reset(pes_27_reset),
    .io_cfg_en(pes_27_io_cfg_en),
    .io_cfg_addr(pes_27_io_cfg_addr),
    .io_cfg_data(pes_27_io_cfg_data),
    .io_en(pes_27_io_en),
    .io_in_0(pes_27_io_in_0),
    .io_in_1(pes_27_io_in_1),
    .io_in_2(pes_27_io_in_2),
    .io_in_3(pes_27_io_in_3),
    .io_in_4(pes_27_io_in_4),
    .io_in_5(pes_27_io_in_5),
    .io_in_6(pes_27_io_in_6),
    .io_in_7(pes_27_io_in_7),
    .io_out_0(pes_27_io_out_0)
  );
  GPE_28 pes_28 ( // @[CGRA.scala 200:20]
    .clock(pes_28_clock),
    .reset(pes_28_reset),
    .io_cfg_en(pes_28_io_cfg_en),
    .io_cfg_addr(pes_28_io_cfg_addr),
    .io_cfg_data(pes_28_io_cfg_data),
    .io_en(pes_28_io_en),
    .io_in_0(pes_28_io_in_0),
    .io_in_1(pes_28_io_in_1),
    .io_in_2(pes_28_io_in_2),
    .io_in_3(pes_28_io_in_3),
    .io_in_4(pes_28_io_in_4),
    .io_in_5(pes_28_io_in_5),
    .io_in_6(pes_28_io_in_6),
    .io_in_7(pes_28_io_in_7),
    .io_out_0(pes_28_io_out_0)
  );
  GPE_29 pes_29 ( // @[CGRA.scala 200:20]
    .clock(pes_29_clock),
    .reset(pes_29_reset),
    .io_cfg_en(pes_29_io_cfg_en),
    .io_cfg_addr(pes_29_io_cfg_addr),
    .io_cfg_data(pes_29_io_cfg_data),
    .io_en(pes_29_io_en),
    .io_in_0(pes_29_io_in_0),
    .io_in_1(pes_29_io_in_1),
    .io_in_2(pes_29_io_in_2),
    .io_in_3(pes_29_io_in_3),
    .io_in_4(pes_29_io_in_4),
    .io_in_5(pes_29_io_in_5),
    .io_in_6(pes_29_io_in_6),
    .io_in_7(pes_29_io_in_7),
    .io_out_0(pes_29_io_out_0)
  );
  GPE_30 pes_30 ( // @[CGRA.scala 200:20]
    .clock(pes_30_clock),
    .reset(pes_30_reset),
    .io_cfg_en(pes_30_io_cfg_en),
    .io_cfg_addr(pes_30_io_cfg_addr),
    .io_cfg_data(pes_30_io_cfg_data),
    .io_en(pes_30_io_en),
    .io_in_0(pes_30_io_in_0),
    .io_in_1(pes_30_io_in_1),
    .io_in_2(pes_30_io_in_2),
    .io_in_3(pes_30_io_in_3),
    .io_in_4(pes_30_io_in_4),
    .io_in_5(pes_30_io_in_5),
    .io_in_6(pes_30_io_in_6),
    .io_in_7(pes_30_io_in_7),
    .io_out_0(pes_30_io_out_0)
  );
  GPE_31 pes_31 ( // @[CGRA.scala 200:20]
    .clock(pes_31_clock),
    .reset(pes_31_reset),
    .io_cfg_en(pes_31_io_cfg_en),
    .io_cfg_addr(pes_31_io_cfg_addr),
    .io_cfg_data(pes_31_io_cfg_data),
    .io_en(pes_31_io_en),
    .io_in_0(pes_31_io_in_0),
    .io_in_1(pes_31_io_in_1),
    .io_in_2(pes_31_io_in_2),
    .io_in_3(pes_31_io_in_3),
    .io_in_4(pes_31_io_in_4),
    .io_in_5(pes_31_io_in_5),
    .io_in_6(pes_31_io_in_6),
    .io_in_7(pes_31_io_in_7),
    .io_out_0(pes_31_io_out_0)
  );
  GPE_32 pes_32 ( // @[CGRA.scala 200:20]
    .clock(pes_32_clock),
    .reset(pes_32_reset),
    .io_cfg_en(pes_32_io_cfg_en),
    .io_cfg_addr(pes_32_io_cfg_addr),
    .io_cfg_data(pes_32_io_cfg_data),
    .io_en(pes_32_io_en),
    .io_in_0(pes_32_io_in_0),
    .io_in_1(pes_32_io_in_1),
    .io_in_2(pes_32_io_in_2),
    .io_in_3(pes_32_io_in_3),
    .io_in_4(pes_32_io_in_4),
    .io_in_5(pes_32_io_in_5),
    .io_in_6(pes_32_io_in_6),
    .io_in_7(pes_32_io_in_7),
    .io_out_0(pes_32_io_out_0)
  );
  GPE_33 pes_33 ( // @[CGRA.scala 200:20]
    .clock(pes_33_clock),
    .reset(pes_33_reset),
    .io_cfg_en(pes_33_io_cfg_en),
    .io_cfg_addr(pes_33_io_cfg_addr),
    .io_cfg_data(pes_33_io_cfg_data),
    .io_en(pes_33_io_en),
    .io_in_0(pes_33_io_in_0),
    .io_in_1(pes_33_io_in_1),
    .io_in_2(pes_33_io_in_2),
    .io_in_3(pes_33_io_in_3),
    .io_in_4(pes_33_io_in_4),
    .io_in_5(pes_33_io_in_5),
    .io_in_6(pes_33_io_in_6),
    .io_in_7(pes_33_io_in_7),
    .io_out_0(pes_33_io_out_0)
  );
  GPE_34 pes_34 ( // @[CGRA.scala 200:20]
    .clock(pes_34_clock),
    .reset(pes_34_reset),
    .io_cfg_en(pes_34_io_cfg_en),
    .io_cfg_addr(pes_34_io_cfg_addr),
    .io_cfg_data(pes_34_io_cfg_data),
    .io_en(pes_34_io_en),
    .io_in_0(pes_34_io_in_0),
    .io_in_1(pes_34_io_in_1),
    .io_in_2(pes_34_io_in_2),
    .io_in_3(pes_34_io_in_3),
    .io_in_4(pes_34_io_in_4),
    .io_in_5(pes_34_io_in_5),
    .io_in_6(pes_34_io_in_6),
    .io_in_7(pes_34_io_in_7),
    .io_out_0(pes_34_io_out_0)
  );
  GPE_35 pes_35 ( // @[CGRA.scala 200:20]
    .clock(pes_35_clock),
    .reset(pes_35_reset),
    .io_cfg_en(pes_35_io_cfg_en),
    .io_cfg_addr(pes_35_io_cfg_addr),
    .io_cfg_data(pes_35_io_cfg_data),
    .io_en(pes_35_io_en),
    .io_in_0(pes_35_io_in_0),
    .io_in_1(pes_35_io_in_1),
    .io_in_2(pes_35_io_in_2),
    .io_in_3(pes_35_io_in_3),
    .io_in_4(pes_35_io_in_4),
    .io_in_5(pes_35_io_in_5),
    .io_in_6(pes_35_io_in_6),
    .io_in_7(pes_35_io_in_7),
    .io_out_0(pes_35_io_out_0)
  );
  GPE_36 pes_36 ( // @[CGRA.scala 200:20]
    .clock(pes_36_clock),
    .reset(pes_36_reset),
    .io_cfg_en(pes_36_io_cfg_en),
    .io_cfg_addr(pes_36_io_cfg_addr),
    .io_cfg_data(pes_36_io_cfg_data),
    .io_en(pes_36_io_en),
    .io_in_0(pes_36_io_in_0),
    .io_in_1(pes_36_io_in_1),
    .io_in_2(pes_36_io_in_2),
    .io_in_3(pes_36_io_in_3),
    .io_in_4(pes_36_io_in_4),
    .io_in_5(pes_36_io_in_5),
    .io_in_6(pes_36_io_in_6),
    .io_in_7(pes_36_io_in_7),
    .io_out_0(pes_36_io_out_0)
  );
  GPE_37 pes_37 ( // @[CGRA.scala 200:20]
    .clock(pes_37_clock),
    .reset(pes_37_reset),
    .io_cfg_en(pes_37_io_cfg_en),
    .io_cfg_addr(pes_37_io_cfg_addr),
    .io_cfg_data(pes_37_io_cfg_data),
    .io_en(pes_37_io_en),
    .io_in_0(pes_37_io_in_0),
    .io_in_1(pes_37_io_in_1),
    .io_in_2(pes_37_io_in_2),
    .io_in_3(pes_37_io_in_3),
    .io_in_4(pes_37_io_in_4),
    .io_in_5(pes_37_io_in_5),
    .io_in_6(pes_37_io_in_6),
    .io_in_7(pes_37_io_in_7),
    .io_out_0(pes_37_io_out_0)
  );
  GPE_38 pes_38 ( // @[CGRA.scala 200:20]
    .clock(pes_38_clock),
    .reset(pes_38_reset),
    .io_cfg_en(pes_38_io_cfg_en),
    .io_cfg_addr(pes_38_io_cfg_addr),
    .io_cfg_data(pes_38_io_cfg_data),
    .io_en(pes_38_io_en),
    .io_in_0(pes_38_io_in_0),
    .io_in_1(pes_38_io_in_1),
    .io_in_2(pes_38_io_in_2),
    .io_in_3(pes_38_io_in_3),
    .io_in_4(pes_38_io_in_4),
    .io_in_5(pes_38_io_in_5),
    .io_in_6(pes_38_io_in_6),
    .io_in_7(pes_38_io_in_7),
    .io_out_0(pes_38_io_out_0)
  );
  GPE_39 pes_39 ( // @[CGRA.scala 200:20]
    .clock(pes_39_clock),
    .reset(pes_39_reset),
    .io_cfg_en(pes_39_io_cfg_en),
    .io_cfg_addr(pes_39_io_cfg_addr),
    .io_cfg_data(pes_39_io_cfg_data),
    .io_en(pes_39_io_en),
    .io_in_0(pes_39_io_in_0),
    .io_in_1(pes_39_io_in_1),
    .io_in_2(pes_39_io_in_2),
    .io_in_3(pes_39_io_in_3),
    .io_in_4(pes_39_io_in_4),
    .io_in_5(pes_39_io_in_5),
    .io_in_6(pes_39_io_in_6),
    .io_in_7(pes_39_io_in_7),
    .io_out_0(pes_39_io_out_0)
  );
  GPE_40 pes_40 ( // @[CGRA.scala 200:20]
    .clock(pes_40_clock),
    .reset(pes_40_reset),
    .io_cfg_en(pes_40_io_cfg_en),
    .io_cfg_addr(pes_40_io_cfg_addr),
    .io_cfg_data(pes_40_io_cfg_data),
    .io_en(pes_40_io_en),
    .io_in_0(pes_40_io_in_0),
    .io_in_1(pes_40_io_in_1),
    .io_in_2(pes_40_io_in_2),
    .io_in_3(pes_40_io_in_3),
    .io_in_4(pes_40_io_in_4),
    .io_in_5(pes_40_io_in_5),
    .io_in_6(pes_40_io_in_6),
    .io_in_7(pes_40_io_in_7),
    .io_out_0(pes_40_io_out_0)
  );
  GPE_41 pes_41 ( // @[CGRA.scala 200:20]
    .clock(pes_41_clock),
    .reset(pes_41_reset),
    .io_cfg_en(pes_41_io_cfg_en),
    .io_cfg_addr(pes_41_io_cfg_addr),
    .io_cfg_data(pes_41_io_cfg_data),
    .io_en(pes_41_io_en),
    .io_in_0(pes_41_io_in_0),
    .io_in_1(pes_41_io_in_1),
    .io_in_2(pes_41_io_in_2),
    .io_in_3(pes_41_io_in_3),
    .io_in_4(pes_41_io_in_4),
    .io_in_5(pes_41_io_in_5),
    .io_in_6(pes_41_io_in_6),
    .io_in_7(pes_41_io_in_7),
    .io_out_0(pes_41_io_out_0)
  );
  GPE_42 pes_42 ( // @[CGRA.scala 200:20]
    .clock(pes_42_clock),
    .reset(pes_42_reset),
    .io_cfg_en(pes_42_io_cfg_en),
    .io_cfg_addr(pes_42_io_cfg_addr),
    .io_cfg_data(pes_42_io_cfg_data),
    .io_en(pes_42_io_en),
    .io_in_0(pes_42_io_in_0),
    .io_in_1(pes_42_io_in_1),
    .io_in_2(pes_42_io_in_2),
    .io_in_3(pes_42_io_in_3),
    .io_in_4(pes_42_io_in_4),
    .io_in_5(pes_42_io_in_5),
    .io_in_6(pes_42_io_in_6),
    .io_in_7(pes_42_io_in_7),
    .io_out_0(pes_42_io_out_0)
  );
  GPE_43 pes_43 ( // @[CGRA.scala 200:20]
    .clock(pes_43_clock),
    .reset(pes_43_reset),
    .io_cfg_en(pes_43_io_cfg_en),
    .io_cfg_addr(pes_43_io_cfg_addr),
    .io_cfg_data(pes_43_io_cfg_data),
    .io_en(pes_43_io_en),
    .io_in_0(pes_43_io_in_0),
    .io_in_1(pes_43_io_in_1),
    .io_in_2(pes_43_io_in_2),
    .io_in_3(pes_43_io_in_3),
    .io_in_4(pes_43_io_in_4),
    .io_in_5(pes_43_io_in_5),
    .io_in_6(pes_43_io_in_6),
    .io_in_7(pes_43_io_in_7),
    .io_out_0(pes_43_io_out_0)
  );
  GPE_44 pes_44 ( // @[CGRA.scala 200:20]
    .clock(pes_44_clock),
    .reset(pes_44_reset),
    .io_cfg_en(pes_44_io_cfg_en),
    .io_cfg_addr(pes_44_io_cfg_addr),
    .io_cfg_data(pes_44_io_cfg_data),
    .io_en(pes_44_io_en),
    .io_in_0(pes_44_io_in_0),
    .io_in_1(pes_44_io_in_1),
    .io_in_2(pes_44_io_in_2),
    .io_in_3(pes_44_io_in_3),
    .io_in_4(pes_44_io_in_4),
    .io_in_5(pes_44_io_in_5),
    .io_in_6(pes_44_io_in_6),
    .io_in_7(pes_44_io_in_7),
    .io_out_0(pes_44_io_out_0)
  );
  GPE_45 pes_45 ( // @[CGRA.scala 200:20]
    .clock(pes_45_clock),
    .reset(pes_45_reset),
    .io_cfg_en(pes_45_io_cfg_en),
    .io_cfg_addr(pes_45_io_cfg_addr),
    .io_cfg_data(pes_45_io_cfg_data),
    .io_en(pes_45_io_en),
    .io_in_0(pes_45_io_in_0),
    .io_in_1(pes_45_io_in_1),
    .io_in_2(pes_45_io_in_2),
    .io_in_3(pes_45_io_in_3),
    .io_in_4(pes_45_io_in_4),
    .io_in_5(pes_45_io_in_5),
    .io_in_6(pes_45_io_in_6),
    .io_in_7(pes_45_io_in_7),
    .io_out_0(pes_45_io_out_0)
  );
  GPE_46 pes_46 ( // @[CGRA.scala 200:20]
    .clock(pes_46_clock),
    .reset(pes_46_reset),
    .io_cfg_en(pes_46_io_cfg_en),
    .io_cfg_addr(pes_46_io_cfg_addr),
    .io_cfg_data(pes_46_io_cfg_data),
    .io_en(pes_46_io_en),
    .io_in_0(pes_46_io_in_0),
    .io_in_1(pes_46_io_in_1),
    .io_in_2(pes_46_io_in_2),
    .io_in_3(pes_46_io_in_3),
    .io_in_4(pes_46_io_in_4),
    .io_in_5(pes_46_io_in_5),
    .io_in_6(pes_46_io_in_6),
    .io_in_7(pes_46_io_in_7),
    .io_out_0(pes_46_io_out_0)
  );
  GPE_47 pes_47 ( // @[CGRA.scala 200:20]
    .clock(pes_47_clock),
    .reset(pes_47_reset),
    .io_cfg_en(pes_47_io_cfg_en),
    .io_cfg_addr(pes_47_io_cfg_addr),
    .io_cfg_data(pes_47_io_cfg_data),
    .io_en(pes_47_io_en),
    .io_in_0(pes_47_io_in_0),
    .io_in_1(pes_47_io_in_1),
    .io_in_2(pes_47_io_in_2),
    .io_in_3(pes_47_io_in_3),
    .io_in_4(pes_47_io_in_4),
    .io_in_5(pes_47_io_in_5),
    .io_in_6(pes_47_io_in_6),
    .io_in_7(pes_47_io_in_7),
    .io_out_0(pes_47_io_out_0)
  );
  GPE_48 pes_48 ( // @[CGRA.scala 200:20]
    .clock(pes_48_clock),
    .reset(pes_48_reset),
    .io_cfg_en(pes_48_io_cfg_en),
    .io_cfg_addr(pes_48_io_cfg_addr),
    .io_cfg_data(pes_48_io_cfg_data),
    .io_en(pes_48_io_en),
    .io_in_0(pes_48_io_in_0),
    .io_in_1(pes_48_io_in_1),
    .io_in_2(pes_48_io_in_2),
    .io_in_3(pes_48_io_in_3),
    .io_in_4(pes_48_io_in_4),
    .io_in_5(pes_48_io_in_5),
    .io_in_6(pes_48_io_in_6),
    .io_in_7(pes_48_io_in_7),
    .io_out_0(pes_48_io_out_0)
  );
  GPE_49 pes_49 ( // @[CGRA.scala 200:20]
    .clock(pes_49_clock),
    .reset(pes_49_reset),
    .io_cfg_en(pes_49_io_cfg_en),
    .io_cfg_addr(pes_49_io_cfg_addr),
    .io_cfg_data(pes_49_io_cfg_data),
    .io_en(pes_49_io_en),
    .io_in_0(pes_49_io_in_0),
    .io_in_1(pes_49_io_in_1),
    .io_in_2(pes_49_io_in_2),
    .io_in_3(pes_49_io_in_3),
    .io_in_4(pes_49_io_in_4),
    .io_in_5(pes_49_io_in_5),
    .io_in_6(pes_49_io_in_6),
    .io_in_7(pes_49_io_in_7),
    .io_out_0(pes_49_io_out_0)
  );
  GPE_50 pes_50 ( // @[CGRA.scala 200:20]
    .clock(pes_50_clock),
    .reset(pes_50_reset),
    .io_cfg_en(pes_50_io_cfg_en),
    .io_cfg_addr(pes_50_io_cfg_addr),
    .io_cfg_data(pes_50_io_cfg_data),
    .io_en(pes_50_io_en),
    .io_in_0(pes_50_io_in_0),
    .io_in_1(pes_50_io_in_1),
    .io_in_2(pes_50_io_in_2),
    .io_in_3(pes_50_io_in_3),
    .io_in_4(pes_50_io_in_4),
    .io_in_5(pes_50_io_in_5),
    .io_in_6(pes_50_io_in_6),
    .io_in_7(pes_50_io_in_7),
    .io_out_0(pes_50_io_out_0)
  );
  GPE_51 pes_51 ( // @[CGRA.scala 200:20]
    .clock(pes_51_clock),
    .reset(pes_51_reset),
    .io_cfg_en(pes_51_io_cfg_en),
    .io_cfg_addr(pes_51_io_cfg_addr),
    .io_cfg_data(pes_51_io_cfg_data),
    .io_en(pes_51_io_en),
    .io_in_0(pes_51_io_in_0),
    .io_in_1(pes_51_io_in_1),
    .io_in_2(pes_51_io_in_2),
    .io_in_3(pes_51_io_in_3),
    .io_in_4(pes_51_io_in_4),
    .io_in_5(pes_51_io_in_5),
    .io_in_6(pes_51_io_in_6),
    .io_in_7(pes_51_io_in_7),
    .io_out_0(pes_51_io_out_0)
  );
  GPE_52 pes_52 ( // @[CGRA.scala 200:20]
    .clock(pes_52_clock),
    .reset(pes_52_reset),
    .io_cfg_en(pes_52_io_cfg_en),
    .io_cfg_addr(pes_52_io_cfg_addr),
    .io_cfg_data(pes_52_io_cfg_data),
    .io_en(pes_52_io_en),
    .io_in_0(pes_52_io_in_0),
    .io_in_1(pes_52_io_in_1),
    .io_in_2(pes_52_io_in_2),
    .io_in_3(pes_52_io_in_3),
    .io_in_4(pes_52_io_in_4),
    .io_in_5(pes_52_io_in_5),
    .io_in_6(pes_52_io_in_6),
    .io_in_7(pes_52_io_in_7),
    .io_out_0(pes_52_io_out_0)
  );
  GPE_53 pes_53 ( // @[CGRA.scala 200:20]
    .clock(pes_53_clock),
    .reset(pes_53_reset),
    .io_cfg_en(pes_53_io_cfg_en),
    .io_cfg_addr(pes_53_io_cfg_addr),
    .io_cfg_data(pes_53_io_cfg_data),
    .io_en(pes_53_io_en),
    .io_in_0(pes_53_io_in_0),
    .io_in_1(pes_53_io_in_1),
    .io_in_2(pes_53_io_in_2),
    .io_in_3(pes_53_io_in_3),
    .io_in_4(pes_53_io_in_4),
    .io_in_5(pes_53_io_in_5),
    .io_in_6(pes_53_io_in_6),
    .io_in_7(pes_53_io_in_7),
    .io_out_0(pes_53_io_out_0)
  );
  GPE_54 pes_54 ( // @[CGRA.scala 200:20]
    .clock(pes_54_clock),
    .reset(pes_54_reset),
    .io_cfg_en(pes_54_io_cfg_en),
    .io_cfg_addr(pes_54_io_cfg_addr),
    .io_cfg_data(pes_54_io_cfg_data),
    .io_en(pes_54_io_en),
    .io_in_0(pes_54_io_in_0),
    .io_in_1(pes_54_io_in_1),
    .io_in_2(pes_54_io_in_2),
    .io_in_3(pes_54_io_in_3),
    .io_in_4(pes_54_io_in_4),
    .io_in_5(pes_54_io_in_5),
    .io_in_6(pes_54_io_in_6),
    .io_in_7(pes_54_io_in_7),
    .io_out_0(pes_54_io_out_0)
  );
  GPE_55 pes_55 ( // @[CGRA.scala 200:20]
    .clock(pes_55_clock),
    .reset(pes_55_reset),
    .io_cfg_en(pes_55_io_cfg_en),
    .io_cfg_addr(pes_55_io_cfg_addr),
    .io_cfg_data(pes_55_io_cfg_data),
    .io_en(pes_55_io_en),
    .io_in_0(pes_55_io_in_0),
    .io_in_1(pes_55_io_in_1),
    .io_in_2(pes_55_io_in_2),
    .io_in_3(pes_55_io_in_3),
    .io_in_4(pes_55_io_in_4),
    .io_in_5(pes_55_io_in_5),
    .io_in_6(pes_55_io_in_6),
    .io_in_7(pes_55_io_in_7),
    .io_out_0(pes_55_io_out_0)
  );
  GPE_56 pes_56 ( // @[CGRA.scala 200:20]
    .clock(pes_56_clock),
    .reset(pes_56_reset),
    .io_cfg_en(pes_56_io_cfg_en),
    .io_cfg_addr(pes_56_io_cfg_addr),
    .io_cfg_data(pes_56_io_cfg_data),
    .io_en(pes_56_io_en),
    .io_in_0(pes_56_io_in_0),
    .io_in_1(pes_56_io_in_1),
    .io_in_2(pes_56_io_in_2),
    .io_in_3(pes_56_io_in_3),
    .io_in_4(pes_56_io_in_4),
    .io_in_5(pes_56_io_in_5),
    .io_in_6(pes_56_io_in_6),
    .io_in_7(pes_56_io_in_7),
    .io_out_0(pes_56_io_out_0)
  );
  GPE_57 pes_57 ( // @[CGRA.scala 200:20]
    .clock(pes_57_clock),
    .reset(pes_57_reset),
    .io_cfg_en(pes_57_io_cfg_en),
    .io_cfg_addr(pes_57_io_cfg_addr),
    .io_cfg_data(pes_57_io_cfg_data),
    .io_en(pes_57_io_en),
    .io_in_0(pes_57_io_in_0),
    .io_in_1(pes_57_io_in_1),
    .io_in_2(pes_57_io_in_2),
    .io_in_3(pes_57_io_in_3),
    .io_in_4(pes_57_io_in_4),
    .io_in_5(pes_57_io_in_5),
    .io_in_6(pes_57_io_in_6),
    .io_in_7(pes_57_io_in_7),
    .io_out_0(pes_57_io_out_0)
  );
  GPE_58 pes_58 ( // @[CGRA.scala 200:20]
    .clock(pes_58_clock),
    .reset(pes_58_reset),
    .io_cfg_en(pes_58_io_cfg_en),
    .io_cfg_addr(pes_58_io_cfg_addr),
    .io_cfg_data(pes_58_io_cfg_data),
    .io_en(pes_58_io_en),
    .io_in_0(pes_58_io_in_0),
    .io_in_1(pes_58_io_in_1),
    .io_in_2(pes_58_io_in_2),
    .io_in_3(pes_58_io_in_3),
    .io_in_4(pes_58_io_in_4),
    .io_in_5(pes_58_io_in_5),
    .io_in_6(pes_58_io_in_6),
    .io_in_7(pes_58_io_in_7),
    .io_out_0(pes_58_io_out_0)
  );
  GPE_59 pes_59 ( // @[CGRA.scala 200:20]
    .clock(pes_59_clock),
    .reset(pes_59_reset),
    .io_cfg_en(pes_59_io_cfg_en),
    .io_cfg_addr(pes_59_io_cfg_addr),
    .io_cfg_data(pes_59_io_cfg_data),
    .io_en(pes_59_io_en),
    .io_in_0(pes_59_io_in_0),
    .io_in_1(pes_59_io_in_1),
    .io_in_2(pes_59_io_in_2),
    .io_in_3(pes_59_io_in_3),
    .io_in_4(pes_59_io_in_4),
    .io_in_5(pes_59_io_in_5),
    .io_in_6(pes_59_io_in_6),
    .io_in_7(pes_59_io_in_7),
    .io_out_0(pes_59_io_out_0)
  );
  GPE_60 pes_60 ( // @[CGRA.scala 200:20]
    .clock(pes_60_clock),
    .reset(pes_60_reset),
    .io_cfg_en(pes_60_io_cfg_en),
    .io_cfg_addr(pes_60_io_cfg_addr),
    .io_cfg_data(pes_60_io_cfg_data),
    .io_en(pes_60_io_en),
    .io_in_0(pes_60_io_in_0),
    .io_in_1(pes_60_io_in_1),
    .io_in_2(pes_60_io_in_2),
    .io_in_3(pes_60_io_in_3),
    .io_in_4(pes_60_io_in_4),
    .io_in_5(pes_60_io_in_5),
    .io_in_6(pes_60_io_in_6),
    .io_in_7(pes_60_io_in_7),
    .io_out_0(pes_60_io_out_0)
  );
  GPE_61 pes_61 ( // @[CGRA.scala 200:20]
    .clock(pes_61_clock),
    .reset(pes_61_reset),
    .io_cfg_en(pes_61_io_cfg_en),
    .io_cfg_addr(pes_61_io_cfg_addr),
    .io_cfg_data(pes_61_io_cfg_data),
    .io_en(pes_61_io_en),
    .io_in_0(pes_61_io_in_0),
    .io_in_1(pes_61_io_in_1),
    .io_in_2(pes_61_io_in_2),
    .io_in_3(pes_61_io_in_3),
    .io_in_4(pes_61_io_in_4),
    .io_in_5(pes_61_io_in_5),
    .io_in_6(pes_61_io_in_6),
    .io_in_7(pes_61_io_in_7),
    .io_out_0(pes_61_io_out_0)
  );
  GPE_62 pes_62 ( // @[CGRA.scala 200:20]
    .clock(pes_62_clock),
    .reset(pes_62_reset),
    .io_cfg_en(pes_62_io_cfg_en),
    .io_cfg_addr(pes_62_io_cfg_addr),
    .io_cfg_data(pes_62_io_cfg_data),
    .io_en(pes_62_io_en),
    .io_in_0(pes_62_io_in_0),
    .io_in_1(pes_62_io_in_1),
    .io_in_2(pes_62_io_in_2),
    .io_in_3(pes_62_io_in_3),
    .io_in_4(pes_62_io_in_4),
    .io_in_5(pes_62_io_in_5),
    .io_in_6(pes_62_io_in_6),
    .io_in_7(pes_62_io_in_7),
    .io_out_0(pes_62_io_out_0)
  );
  GPE_63 pes_63 ( // @[CGRA.scala 200:20]
    .clock(pes_63_clock),
    .reset(pes_63_reset),
    .io_cfg_en(pes_63_io_cfg_en),
    .io_cfg_addr(pes_63_io_cfg_addr),
    .io_cfg_data(pes_63_io_cfg_data),
    .io_en(pes_63_io_en),
    .io_in_0(pes_63_io_in_0),
    .io_in_1(pes_63_io_in_1),
    .io_in_2(pes_63_io_in_2),
    .io_in_3(pes_63_io_in_3),
    .io_in_4(pes_63_io_in_4),
    .io_in_5(pes_63_io_in_5),
    .io_in_6(pes_63_io_in_6),
    .io_in_7(pes_63_io_in_7),
    .io_out_0(pes_63_io_out_0)
  );
  GIB gibs_0 ( // @[CGRA.scala 273:21]
    .clock(gibs_0_clock),
    .reset(gibs_0_reset),
    .io_cfg_en(gibs_0_io_cfg_en),
    .io_cfg_addr(gibs_0_io_cfg_addr),
    .io_cfg_data(gibs_0_io_cfg_data),
    .io_ipinNE_0(gibs_0_io_ipinNE_0),
    .io_opinNE_0(gibs_0_io_opinNE_0),
    .io_ipinSE_0(gibs_0_io_ipinSE_0),
    .io_ipinSE_1(gibs_0_io_ipinSE_1),
    .io_opinSE_0(gibs_0_io_opinSE_0),
    .io_itrackE_0(gibs_0_io_itrackE_0),
    .io_otrackE_0(gibs_0_io_otrackE_0),
    .io_itrackS_0(gibs_0_io_itrackS_0),
    .io_otrackS_0(gibs_0_io_otrackS_0)
  );
  GIB_1 gibs_1 ( // @[CGRA.scala 273:21]
    .clock(gibs_1_clock),
    .reset(gibs_1_reset),
    .io_cfg_en(gibs_1_io_cfg_en),
    .io_cfg_addr(gibs_1_io_cfg_addr),
    .io_cfg_data(gibs_1_io_cfg_data),
    .io_ipinNW_0(gibs_1_io_ipinNW_0),
    .io_opinNW_0(gibs_1_io_opinNW_0),
    .io_ipinNE_0(gibs_1_io_ipinNE_0),
    .io_opinNE_0(gibs_1_io_opinNE_0),
    .io_ipinSE_0(gibs_1_io_ipinSE_0),
    .io_ipinSE_1(gibs_1_io_ipinSE_1),
    .io_opinSE_0(gibs_1_io_opinSE_0),
    .io_ipinSW_0(gibs_1_io_ipinSW_0),
    .io_ipinSW_1(gibs_1_io_ipinSW_1),
    .io_opinSW_0(gibs_1_io_opinSW_0),
    .io_itrackW_0(gibs_1_io_itrackW_0),
    .io_otrackW_0(gibs_1_io_otrackW_0),
    .io_itrackE_0(gibs_1_io_itrackE_0),
    .io_otrackE_0(gibs_1_io_otrackE_0),
    .io_itrackS_0(gibs_1_io_itrackS_0),
    .io_otrackS_0(gibs_1_io_otrackS_0)
  );
  GIB_2 gibs_2 ( // @[CGRA.scala 273:21]
    .clock(gibs_2_clock),
    .reset(gibs_2_reset),
    .io_cfg_en(gibs_2_io_cfg_en),
    .io_cfg_addr(gibs_2_io_cfg_addr),
    .io_cfg_data(gibs_2_io_cfg_data),
    .io_ipinNW_0(gibs_2_io_ipinNW_0),
    .io_opinNW_0(gibs_2_io_opinNW_0),
    .io_ipinNE_0(gibs_2_io_ipinNE_0),
    .io_opinNE_0(gibs_2_io_opinNE_0),
    .io_ipinSE_0(gibs_2_io_ipinSE_0),
    .io_ipinSE_1(gibs_2_io_ipinSE_1),
    .io_opinSE_0(gibs_2_io_opinSE_0),
    .io_ipinSW_0(gibs_2_io_ipinSW_0),
    .io_ipinSW_1(gibs_2_io_ipinSW_1),
    .io_opinSW_0(gibs_2_io_opinSW_0),
    .io_itrackW_0(gibs_2_io_itrackW_0),
    .io_otrackW_0(gibs_2_io_otrackW_0),
    .io_itrackE_0(gibs_2_io_itrackE_0),
    .io_otrackE_0(gibs_2_io_otrackE_0),
    .io_itrackS_0(gibs_2_io_itrackS_0),
    .io_otrackS_0(gibs_2_io_otrackS_0)
  );
  GIB_3 gibs_3 ( // @[CGRA.scala 273:21]
    .clock(gibs_3_clock),
    .reset(gibs_3_reset),
    .io_cfg_en(gibs_3_io_cfg_en),
    .io_cfg_addr(gibs_3_io_cfg_addr),
    .io_cfg_data(gibs_3_io_cfg_data),
    .io_ipinNW_0(gibs_3_io_ipinNW_0),
    .io_opinNW_0(gibs_3_io_opinNW_0),
    .io_ipinNE_0(gibs_3_io_ipinNE_0),
    .io_opinNE_0(gibs_3_io_opinNE_0),
    .io_ipinSE_0(gibs_3_io_ipinSE_0),
    .io_ipinSE_1(gibs_3_io_ipinSE_1),
    .io_opinSE_0(gibs_3_io_opinSE_0),
    .io_ipinSW_0(gibs_3_io_ipinSW_0),
    .io_ipinSW_1(gibs_3_io_ipinSW_1),
    .io_opinSW_0(gibs_3_io_opinSW_0),
    .io_itrackW_0(gibs_3_io_itrackW_0),
    .io_otrackW_0(gibs_3_io_otrackW_0),
    .io_itrackE_0(gibs_3_io_itrackE_0),
    .io_otrackE_0(gibs_3_io_otrackE_0),
    .io_itrackS_0(gibs_3_io_itrackS_0),
    .io_otrackS_0(gibs_3_io_otrackS_0)
  );
  GIB_4 gibs_4 ( // @[CGRA.scala 273:21]
    .clock(gibs_4_clock),
    .reset(gibs_4_reset),
    .io_cfg_en(gibs_4_io_cfg_en),
    .io_cfg_addr(gibs_4_io_cfg_addr),
    .io_cfg_data(gibs_4_io_cfg_data),
    .io_ipinNW_0(gibs_4_io_ipinNW_0),
    .io_opinNW_0(gibs_4_io_opinNW_0),
    .io_ipinNE_0(gibs_4_io_ipinNE_0),
    .io_opinNE_0(gibs_4_io_opinNE_0),
    .io_ipinSE_0(gibs_4_io_ipinSE_0),
    .io_ipinSE_1(gibs_4_io_ipinSE_1),
    .io_opinSE_0(gibs_4_io_opinSE_0),
    .io_ipinSW_0(gibs_4_io_ipinSW_0),
    .io_ipinSW_1(gibs_4_io_ipinSW_1),
    .io_opinSW_0(gibs_4_io_opinSW_0),
    .io_itrackW_0(gibs_4_io_itrackW_0),
    .io_otrackW_0(gibs_4_io_otrackW_0),
    .io_itrackE_0(gibs_4_io_itrackE_0),
    .io_otrackE_0(gibs_4_io_otrackE_0),
    .io_itrackS_0(gibs_4_io_itrackS_0),
    .io_otrackS_0(gibs_4_io_otrackS_0)
  );
  GIB_5 gibs_5 ( // @[CGRA.scala 273:21]
    .clock(gibs_5_clock),
    .reset(gibs_5_reset),
    .io_cfg_en(gibs_5_io_cfg_en),
    .io_cfg_addr(gibs_5_io_cfg_addr),
    .io_cfg_data(gibs_5_io_cfg_data),
    .io_ipinNW_0(gibs_5_io_ipinNW_0),
    .io_opinNW_0(gibs_5_io_opinNW_0),
    .io_ipinNE_0(gibs_5_io_ipinNE_0),
    .io_opinNE_0(gibs_5_io_opinNE_0),
    .io_ipinSE_0(gibs_5_io_ipinSE_0),
    .io_ipinSE_1(gibs_5_io_ipinSE_1),
    .io_opinSE_0(gibs_5_io_opinSE_0),
    .io_ipinSW_0(gibs_5_io_ipinSW_0),
    .io_ipinSW_1(gibs_5_io_ipinSW_1),
    .io_opinSW_0(gibs_5_io_opinSW_0),
    .io_itrackW_0(gibs_5_io_itrackW_0),
    .io_otrackW_0(gibs_5_io_otrackW_0),
    .io_itrackE_0(gibs_5_io_itrackE_0),
    .io_otrackE_0(gibs_5_io_otrackE_0),
    .io_itrackS_0(gibs_5_io_itrackS_0),
    .io_otrackS_0(gibs_5_io_otrackS_0)
  );
  GIB_6 gibs_6 ( // @[CGRA.scala 273:21]
    .clock(gibs_6_clock),
    .reset(gibs_6_reset),
    .io_cfg_en(gibs_6_io_cfg_en),
    .io_cfg_addr(gibs_6_io_cfg_addr),
    .io_cfg_data(gibs_6_io_cfg_data),
    .io_ipinNW_0(gibs_6_io_ipinNW_0),
    .io_opinNW_0(gibs_6_io_opinNW_0),
    .io_ipinNE_0(gibs_6_io_ipinNE_0),
    .io_opinNE_0(gibs_6_io_opinNE_0),
    .io_ipinSE_0(gibs_6_io_ipinSE_0),
    .io_ipinSE_1(gibs_6_io_ipinSE_1),
    .io_opinSE_0(gibs_6_io_opinSE_0),
    .io_ipinSW_0(gibs_6_io_ipinSW_0),
    .io_ipinSW_1(gibs_6_io_ipinSW_1),
    .io_opinSW_0(gibs_6_io_opinSW_0),
    .io_itrackW_0(gibs_6_io_itrackW_0),
    .io_otrackW_0(gibs_6_io_otrackW_0),
    .io_itrackE_0(gibs_6_io_itrackE_0),
    .io_otrackE_0(gibs_6_io_otrackE_0),
    .io_itrackS_0(gibs_6_io_itrackS_0),
    .io_otrackS_0(gibs_6_io_otrackS_0)
  );
  GIB_7 gibs_7 ( // @[CGRA.scala 273:21]
    .clock(gibs_7_clock),
    .reset(gibs_7_reset),
    .io_cfg_en(gibs_7_io_cfg_en),
    .io_cfg_addr(gibs_7_io_cfg_addr),
    .io_cfg_data(gibs_7_io_cfg_data),
    .io_ipinNW_0(gibs_7_io_ipinNW_0),
    .io_opinNW_0(gibs_7_io_opinNW_0),
    .io_ipinNE_0(gibs_7_io_ipinNE_0),
    .io_opinNE_0(gibs_7_io_opinNE_0),
    .io_ipinSE_0(gibs_7_io_ipinSE_0),
    .io_ipinSE_1(gibs_7_io_ipinSE_1),
    .io_opinSE_0(gibs_7_io_opinSE_0),
    .io_ipinSW_0(gibs_7_io_ipinSW_0),
    .io_ipinSW_1(gibs_7_io_ipinSW_1),
    .io_opinSW_0(gibs_7_io_opinSW_0),
    .io_itrackW_0(gibs_7_io_itrackW_0),
    .io_otrackW_0(gibs_7_io_otrackW_0),
    .io_itrackE_0(gibs_7_io_itrackE_0),
    .io_otrackE_0(gibs_7_io_otrackE_0),
    .io_itrackS_0(gibs_7_io_itrackS_0),
    .io_otrackS_0(gibs_7_io_otrackS_0)
  );
  GIB_8 gibs_8 ( // @[CGRA.scala 273:21]
    .clock(gibs_8_clock),
    .reset(gibs_8_reset),
    .io_cfg_en(gibs_8_io_cfg_en),
    .io_cfg_addr(gibs_8_io_cfg_addr),
    .io_cfg_data(gibs_8_io_cfg_data),
    .io_ipinNW_0(gibs_8_io_ipinNW_0),
    .io_opinNW_0(gibs_8_io_opinNW_0),
    .io_ipinSW_0(gibs_8_io_ipinSW_0),
    .io_ipinSW_1(gibs_8_io_ipinSW_1),
    .io_opinSW_0(gibs_8_io_opinSW_0),
    .io_itrackW_0(gibs_8_io_itrackW_0),
    .io_otrackW_0(gibs_8_io_otrackW_0),
    .io_itrackS_0(gibs_8_io_itrackS_0),
    .io_otrackS_0(gibs_8_io_otrackS_0)
  );
  GIB_9 gibs_9 ( // @[CGRA.scala 273:21]
    .clock(gibs_9_clock),
    .reset(gibs_9_reset),
    .io_cfg_en(gibs_9_io_cfg_en),
    .io_cfg_addr(gibs_9_io_cfg_addr),
    .io_cfg_data(gibs_9_io_cfg_data),
    .io_ipinNE_0(gibs_9_io_ipinNE_0),
    .io_ipinNE_1(gibs_9_io_ipinNE_1),
    .io_opinNE_0(gibs_9_io_opinNE_0),
    .io_ipinSE_0(gibs_9_io_ipinSE_0),
    .io_ipinSE_1(gibs_9_io_ipinSE_1),
    .io_opinSE_0(gibs_9_io_opinSE_0),
    .io_itrackN_0(gibs_9_io_itrackN_0),
    .io_otrackN_0(gibs_9_io_otrackN_0),
    .io_itrackE_0(gibs_9_io_itrackE_0),
    .io_otrackE_0(gibs_9_io_otrackE_0),
    .io_itrackS_0(gibs_9_io_itrackS_0),
    .io_otrackS_0(gibs_9_io_otrackS_0)
  );
  GIB_10 gibs_10 ( // @[CGRA.scala 273:21]
    .clock(gibs_10_clock),
    .reset(gibs_10_reset),
    .io_cfg_en(gibs_10_io_cfg_en),
    .io_cfg_addr(gibs_10_io_cfg_addr),
    .io_cfg_data(gibs_10_io_cfg_data),
    .io_ipinNW_0(gibs_10_io_ipinNW_0),
    .io_ipinNW_1(gibs_10_io_ipinNW_1),
    .io_opinNW_0(gibs_10_io_opinNW_0),
    .io_ipinNE_0(gibs_10_io_ipinNE_0),
    .io_ipinNE_1(gibs_10_io_ipinNE_1),
    .io_opinNE_0(gibs_10_io_opinNE_0),
    .io_ipinSE_0(gibs_10_io_ipinSE_0),
    .io_ipinSE_1(gibs_10_io_ipinSE_1),
    .io_opinSE_0(gibs_10_io_opinSE_0),
    .io_ipinSW_0(gibs_10_io_ipinSW_0),
    .io_ipinSW_1(gibs_10_io_ipinSW_1),
    .io_opinSW_0(gibs_10_io_opinSW_0),
    .io_itrackW_0(gibs_10_io_itrackW_0),
    .io_otrackW_0(gibs_10_io_otrackW_0),
    .io_itrackN_0(gibs_10_io_itrackN_0),
    .io_otrackN_0(gibs_10_io_otrackN_0),
    .io_itrackE_0(gibs_10_io_itrackE_0),
    .io_otrackE_0(gibs_10_io_otrackE_0),
    .io_itrackS_0(gibs_10_io_itrackS_0),
    .io_otrackS_0(gibs_10_io_otrackS_0)
  );
  GIB_11 gibs_11 ( // @[CGRA.scala 273:21]
    .clock(gibs_11_clock),
    .reset(gibs_11_reset),
    .io_cfg_en(gibs_11_io_cfg_en),
    .io_cfg_addr(gibs_11_io_cfg_addr),
    .io_cfg_data(gibs_11_io_cfg_data),
    .io_ipinNW_0(gibs_11_io_ipinNW_0),
    .io_ipinNW_1(gibs_11_io_ipinNW_1),
    .io_opinNW_0(gibs_11_io_opinNW_0),
    .io_ipinNE_0(gibs_11_io_ipinNE_0),
    .io_ipinNE_1(gibs_11_io_ipinNE_1),
    .io_opinNE_0(gibs_11_io_opinNE_0),
    .io_ipinSE_0(gibs_11_io_ipinSE_0),
    .io_ipinSE_1(gibs_11_io_ipinSE_1),
    .io_opinSE_0(gibs_11_io_opinSE_0),
    .io_ipinSW_0(gibs_11_io_ipinSW_0),
    .io_ipinSW_1(gibs_11_io_ipinSW_1),
    .io_opinSW_0(gibs_11_io_opinSW_0),
    .io_itrackW_0(gibs_11_io_itrackW_0),
    .io_otrackW_0(gibs_11_io_otrackW_0),
    .io_itrackN_0(gibs_11_io_itrackN_0),
    .io_otrackN_0(gibs_11_io_otrackN_0),
    .io_itrackE_0(gibs_11_io_itrackE_0),
    .io_otrackE_0(gibs_11_io_otrackE_0),
    .io_itrackS_0(gibs_11_io_itrackS_0),
    .io_otrackS_0(gibs_11_io_otrackS_0)
  );
  GIB_12 gibs_12 ( // @[CGRA.scala 273:21]
    .clock(gibs_12_clock),
    .reset(gibs_12_reset),
    .io_cfg_en(gibs_12_io_cfg_en),
    .io_cfg_addr(gibs_12_io_cfg_addr),
    .io_cfg_data(gibs_12_io_cfg_data),
    .io_ipinNW_0(gibs_12_io_ipinNW_0),
    .io_ipinNW_1(gibs_12_io_ipinNW_1),
    .io_opinNW_0(gibs_12_io_opinNW_0),
    .io_ipinNE_0(gibs_12_io_ipinNE_0),
    .io_ipinNE_1(gibs_12_io_ipinNE_1),
    .io_opinNE_0(gibs_12_io_opinNE_0),
    .io_ipinSE_0(gibs_12_io_ipinSE_0),
    .io_ipinSE_1(gibs_12_io_ipinSE_1),
    .io_opinSE_0(gibs_12_io_opinSE_0),
    .io_ipinSW_0(gibs_12_io_ipinSW_0),
    .io_ipinSW_1(gibs_12_io_ipinSW_1),
    .io_opinSW_0(gibs_12_io_opinSW_0),
    .io_itrackW_0(gibs_12_io_itrackW_0),
    .io_otrackW_0(gibs_12_io_otrackW_0),
    .io_itrackN_0(gibs_12_io_itrackN_0),
    .io_otrackN_0(gibs_12_io_otrackN_0),
    .io_itrackE_0(gibs_12_io_itrackE_0),
    .io_otrackE_0(gibs_12_io_otrackE_0),
    .io_itrackS_0(gibs_12_io_itrackS_0),
    .io_otrackS_0(gibs_12_io_otrackS_0)
  );
  GIB_13 gibs_13 ( // @[CGRA.scala 273:21]
    .clock(gibs_13_clock),
    .reset(gibs_13_reset),
    .io_cfg_en(gibs_13_io_cfg_en),
    .io_cfg_addr(gibs_13_io_cfg_addr),
    .io_cfg_data(gibs_13_io_cfg_data),
    .io_ipinNW_0(gibs_13_io_ipinNW_0),
    .io_ipinNW_1(gibs_13_io_ipinNW_1),
    .io_opinNW_0(gibs_13_io_opinNW_0),
    .io_ipinNE_0(gibs_13_io_ipinNE_0),
    .io_ipinNE_1(gibs_13_io_ipinNE_1),
    .io_opinNE_0(gibs_13_io_opinNE_0),
    .io_ipinSE_0(gibs_13_io_ipinSE_0),
    .io_ipinSE_1(gibs_13_io_ipinSE_1),
    .io_opinSE_0(gibs_13_io_opinSE_0),
    .io_ipinSW_0(gibs_13_io_ipinSW_0),
    .io_ipinSW_1(gibs_13_io_ipinSW_1),
    .io_opinSW_0(gibs_13_io_opinSW_0),
    .io_itrackW_0(gibs_13_io_itrackW_0),
    .io_otrackW_0(gibs_13_io_otrackW_0),
    .io_itrackN_0(gibs_13_io_itrackN_0),
    .io_otrackN_0(gibs_13_io_otrackN_0),
    .io_itrackE_0(gibs_13_io_itrackE_0),
    .io_otrackE_0(gibs_13_io_otrackE_0),
    .io_itrackS_0(gibs_13_io_itrackS_0),
    .io_otrackS_0(gibs_13_io_otrackS_0)
  );
  GIB_14 gibs_14 ( // @[CGRA.scala 273:21]
    .clock(gibs_14_clock),
    .reset(gibs_14_reset),
    .io_cfg_en(gibs_14_io_cfg_en),
    .io_cfg_addr(gibs_14_io_cfg_addr),
    .io_cfg_data(gibs_14_io_cfg_data),
    .io_ipinNW_0(gibs_14_io_ipinNW_0),
    .io_ipinNW_1(gibs_14_io_ipinNW_1),
    .io_opinNW_0(gibs_14_io_opinNW_0),
    .io_ipinNE_0(gibs_14_io_ipinNE_0),
    .io_ipinNE_1(gibs_14_io_ipinNE_1),
    .io_opinNE_0(gibs_14_io_opinNE_0),
    .io_ipinSE_0(gibs_14_io_ipinSE_0),
    .io_ipinSE_1(gibs_14_io_ipinSE_1),
    .io_opinSE_0(gibs_14_io_opinSE_0),
    .io_ipinSW_0(gibs_14_io_ipinSW_0),
    .io_ipinSW_1(gibs_14_io_ipinSW_1),
    .io_opinSW_0(gibs_14_io_opinSW_0),
    .io_itrackW_0(gibs_14_io_itrackW_0),
    .io_otrackW_0(gibs_14_io_otrackW_0),
    .io_itrackN_0(gibs_14_io_itrackN_0),
    .io_otrackN_0(gibs_14_io_otrackN_0),
    .io_itrackE_0(gibs_14_io_itrackE_0),
    .io_otrackE_0(gibs_14_io_otrackE_0),
    .io_itrackS_0(gibs_14_io_itrackS_0),
    .io_otrackS_0(gibs_14_io_otrackS_0)
  );
  GIB_15 gibs_15 ( // @[CGRA.scala 273:21]
    .clock(gibs_15_clock),
    .reset(gibs_15_reset),
    .io_cfg_en(gibs_15_io_cfg_en),
    .io_cfg_addr(gibs_15_io_cfg_addr),
    .io_cfg_data(gibs_15_io_cfg_data),
    .io_ipinNW_0(gibs_15_io_ipinNW_0),
    .io_ipinNW_1(gibs_15_io_ipinNW_1),
    .io_opinNW_0(gibs_15_io_opinNW_0),
    .io_ipinNE_0(gibs_15_io_ipinNE_0),
    .io_ipinNE_1(gibs_15_io_ipinNE_1),
    .io_opinNE_0(gibs_15_io_opinNE_0),
    .io_ipinSE_0(gibs_15_io_ipinSE_0),
    .io_ipinSE_1(gibs_15_io_ipinSE_1),
    .io_opinSE_0(gibs_15_io_opinSE_0),
    .io_ipinSW_0(gibs_15_io_ipinSW_0),
    .io_ipinSW_1(gibs_15_io_ipinSW_1),
    .io_opinSW_0(gibs_15_io_opinSW_0),
    .io_itrackW_0(gibs_15_io_itrackW_0),
    .io_otrackW_0(gibs_15_io_otrackW_0),
    .io_itrackN_0(gibs_15_io_itrackN_0),
    .io_otrackN_0(gibs_15_io_otrackN_0),
    .io_itrackE_0(gibs_15_io_itrackE_0),
    .io_otrackE_0(gibs_15_io_otrackE_0),
    .io_itrackS_0(gibs_15_io_itrackS_0),
    .io_otrackS_0(gibs_15_io_otrackS_0)
  );
  GIB_16 gibs_16 ( // @[CGRA.scala 273:21]
    .clock(gibs_16_clock),
    .reset(gibs_16_reset),
    .io_cfg_en(gibs_16_io_cfg_en),
    .io_cfg_addr(gibs_16_io_cfg_addr),
    .io_cfg_data(gibs_16_io_cfg_data),
    .io_ipinNW_0(gibs_16_io_ipinNW_0),
    .io_ipinNW_1(gibs_16_io_ipinNW_1),
    .io_opinNW_0(gibs_16_io_opinNW_0),
    .io_ipinNE_0(gibs_16_io_ipinNE_0),
    .io_ipinNE_1(gibs_16_io_ipinNE_1),
    .io_opinNE_0(gibs_16_io_opinNE_0),
    .io_ipinSE_0(gibs_16_io_ipinSE_0),
    .io_ipinSE_1(gibs_16_io_ipinSE_1),
    .io_opinSE_0(gibs_16_io_opinSE_0),
    .io_ipinSW_0(gibs_16_io_ipinSW_0),
    .io_ipinSW_1(gibs_16_io_ipinSW_1),
    .io_opinSW_0(gibs_16_io_opinSW_0),
    .io_itrackW_0(gibs_16_io_itrackW_0),
    .io_otrackW_0(gibs_16_io_otrackW_0),
    .io_itrackN_0(gibs_16_io_itrackN_0),
    .io_otrackN_0(gibs_16_io_otrackN_0),
    .io_itrackE_0(gibs_16_io_itrackE_0),
    .io_otrackE_0(gibs_16_io_otrackE_0),
    .io_itrackS_0(gibs_16_io_itrackS_0),
    .io_otrackS_0(gibs_16_io_otrackS_0)
  );
  GIB_17 gibs_17 ( // @[CGRA.scala 273:21]
    .clock(gibs_17_clock),
    .reset(gibs_17_reset),
    .io_cfg_en(gibs_17_io_cfg_en),
    .io_cfg_addr(gibs_17_io_cfg_addr),
    .io_cfg_data(gibs_17_io_cfg_data),
    .io_ipinNW_0(gibs_17_io_ipinNW_0),
    .io_ipinNW_1(gibs_17_io_ipinNW_1),
    .io_opinNW_0(gibs_17_io_opinNW_0),
    .io_ipinSW_0(gibs_17_io_ipinSW_0),
    .io_ipinSW_1(gibs_17_io_ipinSW_1),
    .io_opinSW_0(gibs_17_io_opinSW_0),
    .io_itrackW_0(gibs_17_io_itrackW_0),
    .io_otrackW_0(gibs_17_io_otrackW_0),
    .io_itrackN_0(gibs_17_io_itrackN_0),
    .io_otrackN_0(gibs_17_io_otrackN_0),
    .io_itrackS_0(gibs_17_io_itrackS_0),
    .io_otrackS_0(gibs_17_io_otrackS_0)
  );
  GIB_18 gibs_18 ( // @[CGRA.scala 273:21]
    .clock(gibs_18_clock),
    .reset(gibs_18_reset),
    .io_cfg_en(gibs_18_io_cfg_en),
    .io_cfg_addr(gibs_18_io_cfg_addr),
    .io_cfg_data(gibs_18_io_cfg_data),
    .io_ipinNE_0(gibs_18_io_ipinNE_0),
    .io_ipinNE_1(gibs_18_io_ipinNE_1),
    .io_opinNE_0(gibs_18_io_opinNE_0),
    .io_ipinSE_0(gibs_18_io_ipinSE_0),
    .io_ipinSE_1(gibs_18_io_ipinSE_1),
    .io_opinSE_0(gibs_18_io_opinSE_0),
    .io_itrackN_0(gibs_18_io_itrackN_0),
    .io_otrackN_0(gibs_18_io_otrackN_0),
    .io_itrackE_0(gibs_18_io_itrackE_0),
    .io_otrackE_0(gibs_18_io_otrackE_0),
    .io_itrackS_0(gibs_18_io_itrackS_0),
    .io_otrackS_0(gibs_18_io_otrackS_0)
  );
  GIB_19 gibs_19 ( // @[CGRA.scala 273:21]
    .clock(gibs_19_clock),
    .reset(gibs_19_reset),
    .io_cfg_en(gibs_19_io_cfg_en),
    .io_cfg_addr(gibs_19_io_cfg_addr),
    .io_cfg_data(gibs_19_io_cfg_data),
    .io_ipinNW_0(gibs_19_io_ipinNW_0),
    .io_ipinNW_1(gibs_19_io_ipinNW_1),
    .io_opinNW_0(gibs_19_io_opinNW_0),
    .io_ipinNE_0(gibs_19_io_ipinNE_0),
    .io_ipinNE_1(gibs_19_io_ipinNE_1),
    .io_opinNE_0(gibs_19_io_opinNE_0),
    .io_ipinSE_0(gibs_19_io_ipinSE_0),
    .io_ipinSE_1(gibs_19_io_ipinSE_1),
    .io_opinSE_0(gibs_19_io_opinSE_0),
    .io_ipinSW_0(gibs_19_io_ipinSW_0),
    .io_ipinSW_1(gibs_19_io_ipinSW_1),
    .io_opinSW_0(gibs_19_io_opinSW_0),
    .io_itrackW_0(gibs_19_io_itrackW_0),
    .io_otrackW_0(gibs_19_io_otrackW_0),
    .io_itrackN_0(gibs_19_io_itrackN_0),
    .io_otrackN_0(gibs_19_io_otrackN_0),
    .io_itrackE_0(gibs_19_io_itrackE_0),
    .io_otrackE_0(gibs_19_io_otrackE_0),
    .io_itrackS_0(gibs_19_io_itrackS_0),
    .io_otrackS_0(gibs_19_io_otrackS_0)
  );
  GIB_20 gibs_20 ( // @[CGRA.scala 273:21]
    .clock(gibs_20_clock),
    .reset(gibs_20_reset),
    .io_cfg_en(gibs_20_io_cfg_en),
    .io_cfg_addr(gibs_20_io_cfg_addr),
    .io_cfg_data(gibs_20_io_cfg_data),
    .io_ipinNW_0(gibs_20_io_ipinNW_0),
    .io_ipinNW_1(gibs_20_io_ipinNW_1),
    .io_opinNW_0(gibs_20_io_opinNW_0),
    .io_ipinNE_0(gibs_20_io_ipinNE_0),
    .io_ipinNE_1(gibs_20_io_ipinNE_1),
    .io_opinNE_0(gibs_20_io_opinNE_0),
    .io_ipinSE_0(gibs_20_io_ipinSE_0),
    .io_ipinSE_1(gibs_20_io_ipinSE_1),
    .io_opinSE_0(gibs_20_io_opinSE_0),
    .io_ipinSW_0(gibs_20_io_ipinSW_0),
    .io_ipinSW_1(gibs_20_io_ipinSW_1),
    .io_opinSW_0(gibs_20_io_opinSW_0),
    .io_itrackW_0(gibs_20_io_itrackW_0),
    .io_otrackW_0(gibs_20_io_otrackW_0),
    .io_itrackN_0(gibs_20_io_itrackN_0),
    .io_otrackN_0(gibs_20_io_otrackN_0),
    .io_itrackE_0(gibs_20_io_itrackE_0),
    .io_otrackE_0(gibs_20_io_otrackE_0),
    .io_itrackS_0(gibs_20_io_itrackS_0),
    .io_otrackS_0(gibs_20_io_otrackS_0)
  );
  GIB_21 gibs_21 ( // @[CGRA.scala 273:21]
    .clock(gibs_21_clock),
    .reset(gibs_21_reset),
    .io_cfg_en(gibs_21_io_cfg_en),
    .io_cfg_addr(gibs_21_io_cfg_addr),
    .io_cfg_data(gibs_21_io_cfg_data),
    .io_ipinNW_0(gibs_21_io_ipinNW_0),
    .io_ipinNW_1(gibs_21_io_ipinNW_1),
    .io_opinNW_0(gibs_21_io_opinNW_0),
    .io_ipinNE_0(gibs_21_io_ipinNE_0),
    .io_ipinNE_1(gibs_21_io_ipinNE_1),
    .io_opinNE_0(gibs_21_io_opinNE_0),
    .io_ipinSE_0(gibs_21_io_ipinSE_0),
    .io_ipinSE_1(gibs_21_io_ipinSE_1),
    .io_opinSE_0(gibs_21_io_opinSE_0),
    .io_ipinSW_0(gibs_21_io_ipinSW_0),
    .io_ipinSW_1(gibs_21_io_ipinSW_1),
    .io_opinSW_0(gibs_21_io_opinSW_0),
    .io_itrackW_0(gibs_21_io_itrackW_0),
    .io_otrackW_0(gibs_21_io_otrackW_0),
    .io_itrackN_0(gibs_21_io_itrackN_0),
    .io_otrackN_0(gibs_21_io_otrackN_0),
    .io_itrackE_0(gibs_21_io_itrackE_0),
    .io_otrackE_0(gibs_21_io_otrackE_0),
    .io_itrackS_0(gibs_21_io_itrackS_0),
    .io_otrackS_0(gibs_21_io_otrackS_0)
  );
  GIB_22 gibs_22 ( // @[CGRA.scala 273:21]
    .clock(gibs_22_clock),
    .reset(gibs_22_reset),
    .io_cfg_en(gibs_22_io_cfg_en),
    .io_cfg_addr(gibs_22_io_cfg_addr),
    .io_cfg_data(gibs_22_io_cfg_data),
    .io_ipinNW_0(gibs_22_io_ipinNW_0),
    .io_ipinNW_1(gibs_22_io_ipinNW_1),
    .io_opinNW_0(gibs_22_io_opinNW_0),
    .io_ipinNE_0(gibs_22_io_ipinNE_0),
    .io_ipinNE_1(gibs_22_io_ipinNE_1),
    .io_opinNE_0(gibs_22_io_opinNE_0),
    .io_ipinSE_0(gibs_22_io_ipinSE_0),
    .io_ipinSE_1(gibs_22_io_ipinSE_1),
    .io_opinSE_0(gibs_22_io_opinSE_0),
    .io_ipinSW_0(gibs_22_io_ipinSW_0),
    .io_ipinSW_1(gibs_22_io_ipinSW_1),
    .io_opinSW_0(gibs_22_io_opinSW_0),
    .io_itrackW_0(gibs_22_io_itrackW_0),
    .io_otrackW_0(gibs_22_io_otrackW_0),
    .io_itrackN_0(gibs_22_io_itrackN_0),
    .io_otrackN_0(gibs_22_io_otrackN_0),
    .io_itrackE_0(gibs_22_io_itrackE_0),
    .io_otrackE_0(gibs_22_io_otrackE_0),
    .io_itrackS_0(gibs_22_io_itrackS_0),
    .io_otrackS_0(gibs_22_io_otrackS_0)
  );
  GIB_23 gibs_23 ( // @[CGRA.scala 273:21]
    .clock(gibs_23_clock),
    .reset(gibs_23_reset),
    .io_cfg_en(gibs_23_io_cfg_en),
    .io_cfg_addr(gibs_23_io_cfg_addr),
    .io_cfg_data(gibs_23_io_cfg_data),
    .io_ipinNW_0(gibs_23_io_ipinNW_0),
    .io_ipinNW_1(gibs_23_io_ipinNW_1),
    .io_opinNW_0(gibs_23_io_opinNW_0),
    .io_ipinNE_0(gibs_23_io_ipinNE_0),
    .io_ipinNE_1(gibs_23_io_ipinNE_1),
    .io_opinNE_0(gibs_23_io_opinNE_0),
    .io_ipinSE_0(gibs_23_io_ipinSE_0),
    .io_ipinSE_1(gibs_23_io_ipinSE_1),
    .io_opinSE_0(gibs_23_io_opinSE_0),
    .io_ipinSW_0(gibs_23_io_ipinSW_0),
    .io_ipinSW_1(gibs_23_io_ipinSW_1),
    .io_opinSW_0(gibs_23_io_opinSW_0),
    .io_itrackW_0(gibs_23_io_itrackW_0),
    .io_otrackW_0(gibs_23_io_otrackW_0),
    .io_itrackN_0(gibs_23_io_itrackN_0),
    .io_otrackN_0(gibs_23_io_otrackN_0),
    .io_itrackE_0(gibs_23_io_itrackE_0),
    .io_otrackE_0(gibs_23_io_otrackE_0),
    .io_itrackS_0(gibs_23_io_itrackS_0),
    .io_otrackS_0(gibs_23_io_otrackS_0)
  );
  GIB_24 gibs_24 ( // @[CGRA.scala 273:21]
    .clock(gibs_24_clock),
    .reset(gibs_24_reset),
    .io_cfg_en(gibs_24_io_cfg_en),
    .io_cfg_addr(gibs_24_io_cfg_addr),
    .io_cfg_data(gibs_24_io_cfg_data),
    .io_ipinNW_0(gibs_24_io_ipinNW_0),
    .io_ipinNW_1(gibs_24_io_ipinNW_1),
    .io_opinNW_0(gibs_24_io_opinNW_0),
    .io_ipinNE_0(gibs_24_io_ipinNE_0),
    .io_ipinNE_1(gibs_24_io_ipinNE_1),
    .io_opinNE_0(gibs_24_io_opinNE_0),
    .io_ipinSE_0(gibs_24_io_ipinSE_0),
    .io_ipinSE_1(gibs_24_io_ipinSE_1),
    .io_opinSE_0(gibs_24_io_opinSE_0),
    .io_ipinSW_0(gibs_24_io_ipinSW_0),
    .io_ipinSW_1(gibs_24_io_ipinSW_1),
    .io_opinSW_0(gibs_24_io_opinSW_0),
    .io_itrackW_0(gibs_24_io_itrackW_0),
    .io_otrackW_0(gibs_24_io_otrackW_0),
    .io_itrackN_0(gibs_24_io_itrackN_0),
    .io_otrackN_0(gibs_24_io_otrackN_0),
    .io_itrackE_0(gibs_24_io_itrackE_0),
    .io_otrackE_0(gibs_24_io_otrackE_0),
    .io_itrackS_0(gibs_24_io_itrackS_0),
    .io_otrackS_0(gibs_24_io_otrackS_0)
  );
  GIB_25 gibs_25 ( // @[CGRA.scala 273:21]
    .clock(gibs_25_clock),
    .reset(gibs_25_reset),
    .io_cfg_en(gibs_25_io_cfg_en),
    .io_cfg_addr(gibs_25_io_cfg_addr),
    .io_cfg_data(gibs_25_io_cfg_data),
    .io_ipinNW_0(gibs_25_io_ipinNW_0),
    .io_ipinNW_1(gibs_25_io_ipinNW_1),
    .io_opinNW_0(gibs_25_io_opinNW_0),
    .io_ipinNE_0(gibs_25_io_ipinNE_0),
    .io_ipinNE_1(gibs_25_io_ipinNE_1),
    .io_opinNE_0(gibs_25_io_opinNE_0),
    .io_ipinSE_0(gibs_25_io_ipinSE_0),
    .io_ipinSE_1(gibs_25_io_ipinSE_1),
    .io_opinSE_0(gibs_25_io_opinSE_0),
    .io_ipinSW_0(gibs_25_io_ipinSW_0),
    .io_ipinSW_1(gibs_25_io_ipinSW_1),
    .io_opinSW_0(gibs_25_io_opinSW_0),
    .io_itrackW_0(gibs_25_io_itrackW_0),
    .io_otrackW_0(gibs_25_io_otrackW_0),
    .io_itrackN_0(gibs_25_io_itrackN_0),
    .io_otrackN_0(gibs_25_io_otrackN_0),
    .io_itrackE_0(gibs_25_io_itrackE_0),
    .io_otrackE_0(gibs_25_io_otrackE_0),
    .io_itrackS_0(gibs_25_io_itrackS_0),
    .io_otrackS_0(gibs_25_io_otrackS_0)
  );
  GIB_26 gibs_26 ( // @[CGRA.scala 273:21]
    .clock(gibs_26_clock),
    .reset(gibs_26_reset),
    .io_cfg_en(gibs_26_io_cfg_en),
    .io_cfg_addr(gibs_26_io_cfg_addr),
    .io_cfg_data(gibs_26_io_cfg_data),
    .io_ipinNW_0(gibs_26_io_ipinNW_0),
    .io_ipinNW_1(gibs_26_io_ipinNW_1),
    .io_opinNW_0(gibs_26_io_opinNW_0),
    .io_ipinSW_0(gibs_26_io_ipinSW_0),
    .io_ipinSW_1(gibs_26_io_ipinSW_1),
    .io_opinSW_0(gibs_26_io_opinSW_0),
    .io_itrackW_0(gibs_26_io_itrackW_0),
    .io_otrackW_0(gibs_26_io_otrackW_0),
    .io_itrackN_0(gibs_26_io_itrackN_0),
    .io_otrackN_0(gibs_26_io_otrackN_0),
    .io_itrackS_0(gibs_26_io_itrackS_0),
    .io_otrackS_0(gibs_26_io_otrackS_0)
  );
  GIB_27 gibs_27 ( // @[CGRA.scala 273:21]
    .clock(gibs_27_clock),
    .reset(gibs_27_reset),
    .io_cfg_en(gibs_27_io_cfg_en),
    .io_cfg_addr(gibs_27_io_cfg_addr),
    .io_cfg_data(gibs_27_io_cfg_data),
    .io_ipinNE_0(gibs_27_io_ipinNE_0),
    .io_ipinNE_1(gibs_27_io_ipinNE_1),
    .io_opinNE_0(gibs_27_io_opinNE_0),
    .io_ipinSE_0(gibs_27_io_ipinSE_0),
    .io_ipinSE_1(gibs_27_io_ipinSE_1),
    .io_opinSE_0(gibs_27_io_opinSE_0),
    .io_itrackN_0(gibs_27_io_itrackN_0),
    .io_otrackN_0(gibs_27_io_otrackN_0),
    .io_itrackE_0(gibs_27_io_itrackE_0),
    .io_otrackE_0(gibs_27_io_otrackE_0),
    .io_itrackS_0(gibs_27_io_itrackS_0),
    .io_otrackS_0(gibs_27_io_otrackS_0)
  );
  GIB_28 gibs_28 ( // @[CGRA.scala 273:21]
    .clock(gibs_28_clock),
    .reset(gibs_28_reset),
    .io_cfg_en(gibs_28_io_cfg_en),
    .io_cfg_addr(gibs_28_io_cfg_addr),
    .io_cfg_data(gibs_28_io_cfg_data),
    .io_ipinNW_0(gibs_28_io_ipinNW_0),
    .io_ipinNW_1(gibs_28_io_ipinNW_1),
    .io_opinNW_0(gibs_28_io_opinNW_0),
    .io_ipinNE_0(gibs_28_io_ipinNE_0),
    .io_ipinNE_1(gibs_28_io_ipinNE_1),
    .io_opinNE_0(gibs_28_io_opinNE_0),
    .io_ipinSE_0(gibs_28_io_ipinSE_0),
    .io_ipinSE_1(gibs_28_io_ipinSE_1),
    .io_opinSE_0(gibs_28_io_opinSE_0),
    .io_ipinSW_0(gibs_28_io_ipinSW_0),
    .io_ipinSW_1(gibs_28_io_ipinSW_1),
    .io_opinSW_0(gibs_28_io_opinSW_0),
    .io_itrackW_0(gibs_28_io_itrackW_0),
    .io_otrackW_0(gibs_28_io_otrackW_0),
    .io_itrackN_0(gibs_28_io_itrackN_0),
    .io_otrackN_0(gibs_28_io_otrackN_0),
    .io_itrackE_0(gibs_28_io_itrackE_0),
    .io_otrackE_0(gibs_28_io_otrackE_0),
    .io_itrackS_0(gibs_28_io_itrackS_0),
    .io_otrackS_0(gibs_28_io_otrackS_0)
  );
  GIB_29 gibs_29 ( // @[CGRA.scala 273:21]
    .clock(gibs_29_clock),
    .reset(gibs_29_reset),
    .io_cfg_en(gibs_29_io_cfg_en),
    .io_cfg_addr(gibs_29_io_cfg_addr),
    .io_cfg_data(gibs_29_io_cfg_data),
    .io_ipinNW_0(gibs_29_io_ipinNW_0),
    .io_ipinNW_1(gibs_29_io_ipinNW_1),
    .io_opinNW_0(gibs_29_io_opinNW_0),
    .io_ipinNE_0(gibs_29_io_ipinNE_0),
    .io_ipinNE_1(gibs_29_io_ipinNE_1),
    .io_opinNE_0(gibs_29_io_opinNE_0),
    .io_ipinSE_0(gibs_29_io_ipinSE_0),
    .io_ipinSE_1(gibs_29_io_ipinSE_1),
    .io_opinSE_0(gibs_29_io_opinSE_0),
    .io_ipinSW_0(gibs_29_io_ipinSW_0),
    .io_ipinSW_1(gibs_29_io_ipinSW_1),
    .io_opinSW_0(gibs_29_io_opinSW_0),
    .io_itrackW_0(gibs_29_io_itrackW_0),
    .io_otrackW_0(gibs_29_io_otrackW_0),
    .io_itrackN_0(gibs_29_io_itrackN_0),
    .io_otrackN_0(gibs_29_io_otrackN_0),
    .io_itrackE_0(gibs_29_io_itrackE_0),
    .io_otrackE_0(gibs_29_io_otrackE_0),
    .io_itrackS_0(gibs_29_io_itrackS_0),
    .io_otrackS_0(gibs_29_io_otrackS_0)
  );
  GIB_30 gibs_30 ( // @[CGRA.scala 273:21]
    .clock(gibs_30_clock),
    .reset(gibs_30_reset),
    .io_cfg_en(gibs_30_io_cfg_en),
    .io_cfg_addr(gibs_30_io_cfg_addr),
    .io_cfg_data(gibs_30_io_cfg_data),
    .io_ipinNW_0(gibs_30_io_ipinNW_0),
    .io_ipinNW_1(gibs_30_io_ipinNW_1),
    .io_opinNW_0(gibs_30_io_opinNW_0),
    .io_ipinNE_0(gibs_30_io_ipinNE_0),
    .io_ipinNE_1(gibs_30_io_ipinNE_1),
    .io_opinNE_0(gibs_30_io_opinNE_0),
    .io_ipinSE_0(gibs_30_io_ipinSE_0),
    .io_ipinSE_1(gibs_30_io_ipinSE_1),
    .io_opinSE_0(gibs_30_io_opinSE_0),
    .io_ipinSW_0(gibs_30_io_ipinSW_0),
    .io_ipinSW_1(gibs_30_io_ipinSW_1),
    .io_opinSW_0(gibs_30_io_opinSW_0),
    .io_itrackW_0(gibs_30_io_itrackW_0),
    .io_otrackW_0(gibs_30_io_otrackW_0),
    .io_itrackN_0(gibs_30_io_itrackN_0),
    .io_otrackN_0(gibs_30_io_otrackN_0),
    .io_itrackE_0(gibs_30_io_itrackE_0),
    .io_otrackE_0(gibs_30_io_otrackE_0),
    .io_itrackS_0(gibs_30_io_itrackS_0),
    .io_otrackS_0(gibs_30_io_otrackS_0)
  );
  GIB_31 gibs_31 ( // @[CGRA.scala 273:21]
    .clock(gibs_31_clock),
    .reset(gibs_31_reset),
    .io_cfg_en(gibs_31_io_cfg_en),
    .io_cfg_addr(gibs_31_io_cfg_addr),
    .io_cfg_data(gibs_31_io_cfg_data),
    .io_ipinNW_0(gibs_31_io_ipinNW_0),
    .io_ipinNW_1(gibs_31_io_ipinNW_1),
    .io_opinNW_0(gibs_31_io_opinNW_0),
    .io_ipinNE_0(gibs_31_io_ipinNE_0),
    .io_ipinNE_1(gibs_31_io_ipinNE_1),
    .io_opinNE_0(gibs_31_io_opinNE_0),
    .io_ipinSE_0(gibs_31_io_ipinSE_0),
    .io_ipinSE_1(gibs_31_io_ipinSE_1),
    .io_opinSE_0(gibs_31_io_opinSE_0),
    .io_ipinSW_0(gibs_31_io_ipinSW_0),
    .io_ipinSW_1(gibs_31_io_ipinSW_1),
    .io_opinSW_0(gibs_31_io_opinSW_0),
    .io_itrackW_0(gibs_31_io_itrackW_0),
    .io_otrackW_0(gibs_31_io_otrackW_0),
    .io_itrackN_0(gibs_31_io_itrackN_0),
    .io_otrackN_0(gibs_31_io_otrackN_0),
    .io_itrackE_0(gibs_31_io_itrackE_0),
    .io_otrackE_0(gibs_31_io_otrackE_0),
    .io_itrackS_0(gibs_31_io_itrackS_0),
    .io_otrackS_0(gibs_31_io_otrackS_0)
  );
  GIB_32 gibs_32 ( // @[CGRA.scala 273:21]
    .clock(gibs_32_clock),
    .reset(gibs_32_reset),
    .io_cfg_en(gibs_32_io_cfg_en),
    .io_cfg_addr(gibs_32_io_cfg_addr),
    .io_cfg_data(gibs_32_io_cfg_data),
    .io_ipinNW_0(gibs_32_io_ipinNW_0),
    .io_ipinNW_1(gibs_32_io_ipinNW_1),
    .io_opinNW_0(gibs_32_io_opinNW_0),
    .io_ipinNE_0(gibs_32_io_ipinNE_0),
    .io_ipinNE_1(gibs_32_io_ipinNE_1),
    .io_opinNE_0(gibs_32_io_opinNE_0),
    .io_ipinSE_0(gibs_32_io_ipinSE_0),
    .io_ipinSE_1(gibs_32_io_ipinSE_1),
    .io_opinSE_0(gibs_32_io_opinSE_0),
    .io_ipinSW_0(gibs_32_io_ipinSW_0),
    .io_ipinSW_1(gibs_32_io_ipinSW_1),
    .io_opinSW_0(gibs_32_io_opinSW_0),
    .io_itrackW_0(gibs_32_io_itrackW_0),
    .io_otrackW_0(gibs_32_io_otrackW_0),
    .io_itrackN_0(gibs_32_io_itrackN_0),
    .io_otrackN_0(gibs_32_io_otrackN_0),
    .io_itrackE_0(gibs_32_io_itrackE_0),
    .io_otrackE_0(gibs_32_io_otrackE_0),
    .io_itrackS_0(gibs_32_io_itrackS_0),
    .io_otrackS_0(gibs_32_io_otrackS_0)
  );
  GIB_33 gibs_33 ( // @[CGRA.scala 273:21]
    .clock(gibs_33_clock),
    .reset(gibs_33_reset),
    .io_cfg_en(gibs_33_io_cfg_en),
    .io_cfg_addr(gibs_33_io_cfg_addr),
    .io_cfg_data(gibs_33_io_cfg_data),
    .io_ipinNW_0(gibs_33_io_ipinNW_0),
    .io_ipinNW_1(gibs_33_io_ipinNW_1),
    .io_opinNW_0(gibs_33_io_opinNW_0),
    .io_ipinNE_0(gibs_33_io_ipinNE_0),
    .io_ipinNE_1(gibs_33_io_ipinNE_1),
    .io_opinNE_0(gibs_33_io_opinNE_0),
    .io_ipinSE_0(gibs_33_io_ipinSE_0),
    .io_ipinSE_1(gibs_33_io_ipinSE_1),
    .io_opinSE_0(gibs_33_io_opinSE_0),
    .io_ipinSW_0(gibs_33_io_ipinSW_0),
    .io_ipinSW_1(gibs_33_io_ipinSW_1),
    .io_opinSW_0(gibs_33_io_opinSW_0),
    .io_itrackW_0(gibs_33_io_itrackW_0),
    .io_otrackW_0(gibs_33_io_otrackW_0),
    .io_itrackN_0(gibs_33_io_itrackN_0),
    .io_otrackN_0(gibs_33_io_otrackN_0),
    .io_itrackE_0(gibs_33_io_itrackE_0),
    .io_otrackE_0(gibs_33_io_otrackE_0),
    .io_itrackS_0(gibs_33_io_itrackS_0),
    .io_otrackS_0(gibs_33_io_otrackS_0)
  );
  GIB_34 gibs_34 ( // @[CGRA.scala 273:21]
    .clock(gibs_34_clock),
    .reset(gibs_34_reset),
    .io_cfg_en(gibs_34_io_cfg_en),
    .io_cfg_addr(gibs_34_io_cfg_addr),
    .io_cfg_data(gibs_34_io_cfg_data),
    .io_ipinNW_0(gibs_34_io_ipinNW_0),
    .io_ipinNW_1(gibs_34_io_ipinNW_1),
    .io_opinNW_0(gibs_34_io_opinNW_0),
    .io_ipinNE_0(gibs_34_io_ipinNE_0),
    .io_ipinNE_1(gibs_34_io_ipinNE_1),
    .io_opinNE_0(gibs_34_io_opinNE_0),
    .io_ipinSE_0(gibs_34_io_ipinSE_0),
    .io_ipinSE_1(gibs_34_io_ipinSE_1),
    .io_opinSE_0(gibs_34_io_opinSE_0),
    .io_ipinSW_0(gibs_34_io_ipinSW_0),
    .io_ipinSW_1(gibs_34_io_ipinSW_1),
    .io_opinSW_0(gibs_34_io_opinSW_0),
    .io_itrackW_0(gibs_34_io_itrackW_0),
    .io_otrackW_0(gibs_34_io_otrackW_0),
    .io_itrackN_0(gibs_34_io_itrackN_0),
    .io_otrackN_0(gibs_34_io_otrackN_0),
    .io_itrackE_0(gibs_34_io_itrackE_0),
    .io_otrackE_0(gibs_34_io_otrackE_0),
    .io_itrackS_0(gibs_34_io_itrackS_0),
    .io_otrackS_0(gibs_34_io_otrackS_0)
  );
  GIB_35 gibs_35 ( // @[CGRA.scala 273:21]
    .clock(gibs_35_clock),
    .reset(gibs_35_reset),
    .io_cfg_en(gibs_35_io_cfg_en),
    .io_cfg_addr(gibs_35_io_cfg_addr),
    .io_cfg_data(gibs_35_io_cfg_data),
    .io_ipinNW_0(gibs_35_io_ipinNW_0),
    .io_ipinNW_1(gibs_35_io_ipinNW_1),
    .io_opinNW_0(gibs_35_io_opinNW_0),
    .io_ipinSW_0(gibs_35_io_ipinSW_0),
    .io_ipinSW_1(gibs_35_io_ipinSW_1),
    .io_opinSW_0(gibs_35_io_opinSW_0),
    .io_itrackW_0(gibs_35_io_itrackW_0),
    .io_otrackW_0(gibs_35_io_otrackW_0),
    .io_itrackN_0(gibs_35_io_itrackN_0),
    .io_otrackN_0(gibs_35_io_otrackN_0),
    .io_itrackS_0(gibs_35_io_itrackS_0),
    .io_otrackS_0(gibs_35_io_otrackS_0)
  );
  GIB_36 gibs_36 ( // @[CGRA.scala 273:21]
    .clock(gibs_36_clock),
    .reset(gibs_36_reset),
    .io_cfg_en(gibs_36_io_cfg_en),
    .io_cfg_addr(gibs_36_io_cfg_addr),
    .io_cfg_data(gibs_36_io_cfg_data),
    .io_ipinNE_0(gibs_36_io_ipinNE_0),
    .io_ipinNE_1(gibs_36_io_ipinNE_1),
    .io_opinNE_0(gibs_36_io_opinNE_0),
    .io_ipinSE_0(gibs_36_io_ipinSE_0),
    .io_ipinSE_1(gibs_36_io_ipinSE_1),
    .io_opinSE_0(gibs_36_io_opinSE_0),
    .io_itrackN_0(gibs_36_io_itrackN_0),
    .io_otrackN_0(gibs_36_io_otrackN_0),
    .io_itrackE_0(gibs_36_io_itrackE_0),
    .io_otrackE_0(gibs_36_io_otrackE_0),
    .io_itrackS_0(gibs_36_io_itrackS_0),
    .io_otrackS_0(gibs_36_io_otrackS_0)
  );
  GIB_37 gibs_37 ( // @[CGRA.scala 273:21]
    .clock(gibs_37_clock),
    .reset(gibs_37_reset),
    .io_cfg_en(gibs_37_io_cfg_en),
    .io_cfg_addr(gibs_37_io_cfg_addr),
    .io_cfg_data(gibs_37_io_cfg_data),
    .io_ipinNW_0(gibs_37_io_ipinNW_0),
    .io_ipinNW_1(gibs_37_io_ipinNW_1),
    .io_opinNW_0(gibs_37_io_opinNW_0),
    .io_ipinNE_0(gibs_37_io_ipinNE_0),
    .io_ipinNE_1(gibs_37_io_ipinNE_1),
    .io_opinNE_0(gibs_37_io_opinNE_0),
    .io_ipinSE_0(gibs_37_io_ipinSE_0),
    .io_ipinSE_1(gibs_37_io_ipinSE_1),
    .io_opinSE_0(gibs_37_io_opinSE_0),
    .io_ipinSW_0(gibs_37_io_ipinSW_0),
    .io_ipinSW_1(gibs_37_io_ipinSW_1),
    .io_opinSW_0(gibs_37_io_opinSW_0),
    .io_itrackW_0(gibs_37_io_itrackW_0),
    .io_otrackW_0(gibs_37_io_otrackW_0),
    .io_itrackN_0(gibs_37_io_itrackN_0),
    .io_otrackN_0(gibs_37_io_otrackN_0),
    .io_itrackE_0(gibs_37_io_itrackE_0),
    .io_otrackE_0(gibs_37_io_otrackE_0),
    .io_itrackS_0(gibs_37_io_itrackS_0),
    .io_otrackS_0(gibs_37_io_otrackS_0)
  );
  GIB_38 gibs_38 ( // @[CGRA.scala 273:21]
    .clock(gibs_38_clock),
    .reset(gibs_38_reset),
    .io_cfg_en(gibs_38_io_cfg_en),
    .io_cfg_addr(gibs_38_io_cfg_addr),
    .io_cfg_data(gibs_38_io_cfg_data),
    .io_ipinNW_0(gibs_38_io_ipinNW_0),
    .io_ipinNW_1(gibs_38_io_ipinNW_1),
    .io_opinNW_0(gibs_38_io_opinNW_0),
    .io_ipinNE_0(gibs_38_io_ipinNE_0),
    .io_ipinNE_1(gibs_38_io_ipinNE_1),
    .io_opinNE_0(gibs_38_io_opinNE_0),
    .io_ipinSE_0(gibs_38_io_ipinSE_0),
    .io_ipinSE_1(gibs_38_io_ipinSE_1),
    .io_opinSE_0(gibs_38_io_opinSE_0),
    .io_ipinSW_0(gibs_38_io_ipinSW_0),
    .io_ipinSW_1(gibs_38_io_ipinSW_1),
    .io_opinSW_0(gibs_38_io_opinSW_0),
    .io_itrackW_0(gibs_38_io_itrackW_0),
    .io_otrackW_0(gibs_38_io_otrackW_0),
    .io_itrackN_0(gibs_38_io_itrackN_0),
    .io_otrackN_0(gibs_38_io_otrackN_0),
    .io_itrackE_0(gibs_38_io_itrackE_0),
    .io_otrackE_0(gibs_38_io_otrackE_0),
    .io_itrackS_0(gibs_38_io_itrackS_0),
    .io_otrackS_0(gibs_38_io_otrackS_0)
  );
  GIB_39 gibs_39 ( // @[CGRA.scala 273:21]
    .clock(gibs_39_clock),
    .reset(gibs_39_reset),
    .io_cfg_en(gibs_39_io_cfg_en),
    .io_cfg_addr(gibs_39_io_cfg_addr),
    .io_cfg_data(gibs_39_io_cfg_data),
    .io_ipinNW_0(gibs_39_io_ipinNW_0),
    .io_ipinNW_1(gibs_39_io_ipinNW_1),
    .io_opinNW_0(gibs_39_io_opinNW_0),
    .io_ipinNE_0(gibs_39_io_ipinNE_0),
    .io_ipinNE_1(gibs_39_io_ipinNE_1),
    .io_opinNE_0(gibs_39_io_opinNE_0),
    .io_ipinSE_0(gibs_39_io_ipinSE_0),
    .io_ipinSE_1(gibs_39_io_ipinSE_1),
    .io_opinSE_0(gibs_39_io_opinSE_0),
    .io_ipinSW_0(gibs_39_io_ipinSW_0),
    .io_ipinSW_1(gibs_39_io_ipinSW_1),
    .io_opinSW_0(gibs_39_io_opinSW_0),
    .io_itrackW_0(gibs_39_io_itrackW_0),
    .io_otrackW_0(gibs_39_io_otrackW_0),
    .io_itrackN_0(gibs_39_io_itrackN_0),
    .io_otrackN_0(gibs_39_io_otrackN_0),
    .io_itrackE_0(gibs_39_io_itrackE_0),
    .io_otrackE_0(gibs_39_io_otrackE_0),
    .io_itrackS_0(gibs_39_io_itrackS_0),
    .io_otrackS_0(gibs_39_io_otrackS_0)
  );
  GIB_40 gibs_40 ( // @[CGRA.scala 273:21]
    .clock(gibs_40_clock),
    .reset(gibs_40_reset),
    .io_cfg_en(gibs_40_io_cfg_en),
    .io_cfg_addr(gibs_40_io_cfg_addr),
    .io_cfg_data(gibs_40_io_cfg_data),
    .io_ipinNW_0(gibs_40_io_ipinNW_0),
    .io_ipinNW_1(gibs_40_io_ipinNW_1),
    .io_opinNW_0(gibs_40_io_opinNW_0),
    .io_ipinNE_0(gibs_40_io_ipinNE_0),
    .io_ipinNE_1(gibs_40_io_ipinNE_1),
    .io_opinNE_0(gibs_40_io_opinNE_0),
    .io_ipinSE_0(gibs_40_io_ipinSE_0),
    .io_ipinSE_1(gibs_40_io_ipinSE_1),
    .io_opinSE_0(gibs_40_io_opinSE_0),
    .io_ipinSW_0(gibs_40_io_ipinSW_0),
    .io_ipinSW_1(gibs_40_io_ipinSW_1),
    .io_opinSW_0(gibs_40_io_opinSW_0),
    .io_itrackW_0(gibs_40_io_itrackW_0),
    .io_otrackW_0(gibs_40_io_otrackW_0),
    .io_itrackN_0(gibs_40_io_itrackN_0),
    .io_otrackN_0(gibs_40_io_otrackN_0),
    .io_itrackE_0(gibs_40_io_itrackE_0),
    .io_otrackE_0(gibs_40_io_otrackE_0),
    .io_itrackS_0(gibs_40_io_itrackS_0),
    .io_otrackS_0(gibs_40_io_otrackS_0)
  );
  GIB_41 gibs_41 ( // @[CGRA.scala 273:21]
    .clock(gibs_41_clock),
    .reset(gibs_41_reset),
    .io_cfg_en(gibs_41_io_cfg_en),
    .io_cfg_addr(gibs_41_io_cfg_addr),
    .io_cfg_data(gibs_41_io_cfg_data),
    .io_ipinNW_0(gibs_41_io_ipinNW_0),
    .io_ipinNW_1(gibs_41_io_ipinNW_1),
    .io_opinNW_0(gibs_41_io_opinNW_0),
    .io_ipinNE_0(gibs_41_io_ipinNE_0),
    .io_ipinNE_1(gibs_41_io_ipinNE_1),
    .io_opinNE_0(gibs_41_io_opinNE_0),
    .io_ipinSE_0(gibs_41_io_ipinSE_0),
    .io_ipinSE_1(gibs_41_io_ipinSE_1),
    .io_opinSE_0(gibs_41_io_opinSE_0),
    .io_ipinSW_0(gibs_41_io_ipinSW_0),
    .io_ipinSW_1(gibs_41_io_ipinSW_1),
    .io_opinSW_0(gibs_41_io_opinSW_0),
    .io_itrackW_0(gibs_41_io_itrackW_0),
    .io_otrackW_0(gibs_41_io_otrackW_0),
    .io_itrackN_0(gibs_41_io_itrackN_0),
    .io_otrackN_0(gibs_41_io_otrackN_0),
    .io_itrackE_0(gibs_41_io_itrackE_0),
    .io_otrackE_0(gibs_41_io_otrackE_0),
    .io_itrackS_0(gibs_41_io_itrackS_0),
    .io_otrackS_0(gibs_41_io_otrackS_0)
  );
  GIB_42 gibs_42 ( // @[CGRA.scala 273:21]
    .clock(gibs_42_clock),
    .reset(gibs_42_reset),
    .io_cfg_en(gibs_42_io_cfg_en),
    .io_cfg_addr(gibs_42_io_cfg_addr),
    .io_cfg_data(gibs_42_io_cfg_data),
    .io_ipinNW_0(gibs_42_io_ipinNW_0),
    .io_ipinNW_1(gibs_42_io_ipinNW_1),
    .io_opinNW_0(gibs_42_io_opinNW_0),
    .io_ipinNE_0(gibs_42_io_ipinNE_0),
    .io_ipinNE_1(gibs_42_io_ipinNE_1),
    .io_opinNE_0(gibs_42_io_opinNE_0),
    .io_ipinSE_0(gibs_42_io_ipinSE_0),
    .io_ipinSE_1(gibs_42_io_ipinSE_1),
    .io_opinSE_0(gibs_42_io_opinSE_0),
    .io_ipinSW_0(gibs_42_io_ipinSW_0),
    .io_ipinSW_1(gibs_42_io_ipinSW_1),
    .io_opinSW_0(gibs_42_io_opinSW_0),
    .io_itrackW_0(gibs_42_io_itrackW_0),
    .io_otrackW_0(gibs_42_io_otrackW_0),
    .io_itrackN_0(gibs_42_io_itrackN_0),
    .io_otrackN_0(gibs_42_io_otrackN_0),
    .io_itrackE_0(gibs_42_io_itrackE_0),
    .io_otrackE_0(gibs_42_io_otrackE_0),
    .io_itrackS_0(gibs_42_io_itrackS_0),
    .io_otrackS_0(gibs_42_io_otrackS_0)
  );
  GIB_43 gibs_43 ( // @[CGRA.scala 273:21]
    .clock(gibs_43_clock),
    .reset(gibs_43_reset),
    .io_cfg_en(gibs_43_io_cfg_en),
    .io_cfg_addr(gibs_43_io_cfg_addr),
    .io_cfg_data(gibs_43_io_cfg_data),
    .io_ipinNW_0(gibs_43_io_ipinNW_0),
    .io_ipinNW_1(gibs_43_io_ipinNW_1),
    .io_opinNW_0(gibs_43_io_opinNW_0),
    .io_ipinNE_0(gibs_43_io_ipinNE_0),
    .io_ipinNE_1(gibs_43_io_ipinNE_1),
    .io_opinNE_0(gibs_43_io_opinNE_0),
    .io_ipinSE_0(gibs_43_io_ipinSE_0),
    .io_ipinSE_1(gibs_43_io_ipinSE_1),
    .io_opinSE_0(gibs_43_io_opinSE_0),
    .io_ipinSW_0(gibs_43_io_ipinSW_0),
    .io_ipinSW_1(gibs_43_io_ipinSW_1),
    .io_opinSW_0(gibs_43_io_opinSW_0),
    .io_itrackW_0(gibs_43_io_itrackW_0),
    .io_otrackW_0(gibs_43_io_otrackW_0),
    .io_itrackN_0(gibs_43_io_itrackN_0),
    .io_otrackN_0(gibs_43_io_otrackN_0),
    .io_itrackE_0(gibs_43_io_itrackE_0),
    .io_otrackE_0(gibs_43_io_otrackE_0),
    .io_itrackS_0(gibs_43_io_itrackS_0),
    .io_otrackS_0(gibs_43_io_otrackS_0)
  );
  GIB_44 gibs_44 ( // @[CGRA.scala 273:21]
    .clock(gibs_44_clock),
    .reset(gibs_44_reset),
    .io_cfg_en(gibs_44_io_cfg_en),
    .io_cfg_addr(gibs_44_io_cfg_addr),
    .io_cfg_data(gibs_44_io_cfg_data),
    .io_ipinNW_0(gibs_44_io_ipinNW_0),
    .io_ipinNW_1(gibs_44_io_ipinNW_1),
    .io_opinNW_0(gibs_44_io_opinNW_0),
    .io_ipinSW_0(gibs_44_io_ipinSW_0),
    .io_ipinSW_1(gibs_44_io_ipinSW_1),
    .io_opinSW_0(gibs_44_io_opinSW_0),
    .io_itrackW_0(gibs_44_io_itrackW_0),
    .io_otrackW_0(gibs_44_io_otrackW_0),
    .io_itrackN_0(gibs_44_io_itrackN_0),
    .io_otrackN_0(gibs_44_io_otrackN_0),
    .io_itrackS_0(gibs_44_io_itrackS_0),
    .io_otrackS_0(gibs_44_io_otrackS_0)
  );
  GIB_45 gibs_45 ( // @[CGRA.scala 273:21]
    .clock(gibs_45_clock),
    .reset(gibs_45_reset),
    .io_cfg_en(gibs_45_io_cfg_en),
    .io_cfg_addr(gibs_45_io_cfg_addr),
    .io_cfg_data(gibs_45_io_cfg_data),
    .io_ipinNE_0(gibs_45_io_ipinNE_0),
    .io_ipinNE_1(gibs_45_io_ipinNE_1),
    .io_opinNE_0(gibs_45_io_opinNE_0),
    .io_ipinSE_0(gibs_45_io_ipinSE_0),
    .io_ipinSE_1(gibs_45_io_ipinSE_1),
    .io_opinSE_0(gibs_45_io_opinSE_0),
    .io_itrackN_0(gibs_45_io_itrackN_0),
    .io_otrackN_0(gibs_45_io_otrackN_0),
    .io_itrackE_0(gibs_45_io_itrackE_0),
    .io_otrackE_0(gibs_45_io_otrackE_0),
    .io_itrackS_0(gibs_45_io_itrackS_0),
    .io_otrackS_0(gibs_45_io_otrackS_0)
  );
  GIB_46 gibs_46 ( // @[CGRA.scala 273:21]
    .clock(gibs_46_clock),
    .reset(gibs_46_reset),
    .io_cfg_en(gibs_46_io_cfg_en),
    .io_cfg_addr(gibs_46_io_cfg_addr),
    .io_cfg_data(gibs_46_io_cfg_data),
    .io_ipinNW_0(gibs_46_io_ipinNW_0),
    .io_ipinNW_1(gibs_46_io_ipinNW_1),
    .io_opinNW_0(gibs_46_io_opinNW_0),
    .io_ipinNE_0(gibs_46_io_ipinNE_0),
    .io_ipinNE_1(gibs_46_io_ipinNE_1),
    .io_opinNE_0(gibs_46_io_opinNE_0),
    .io_ipinSE_0(gibs_46_io_ipinSE_0),
    .io_ipinSE_1(gibs_46_io_ipinSE_1),
    .io_opinSE_0(gibs_46_io_opinSE_0),
    .io_ipinSW_0(gibs_46_io_ipinSW_0),
    .io_ipinSW_1(gibs_46_io_ipinSW_1),
    .io_opinSW_0(gibs_46_io_opinSW_0),
    .io_itrackW_0(gibs_46_io_itrackW_0),
    .io_otrackW_0(gibs_46_io_otrackW_0),
    .io_itrackN_0(gibs_46_io_itrackN_0),
    .io_otrackN_0(gibs_46_io_otrackN_0),
    .io_itrackE_0(gibs_46_io_itrackE_0),
    .io_otrackE_0(gibs_46_io_otrackE_0),
    .io_itrackS_0(gibs_46_io_itrackS_0),
    .io_otrackS_0(gibs_46_io_otrackS_0)
  );
  GIB_47 gibs_47 ( // @[CGRA.scala 273:21]
    .clock(gibs_47_clock),
    .reset(gibs_47_reset),
    .io_cfg_en(gibs_47_io_cfg_en),
    .io_cfg_addr(gibs_47_io_cfg_addr),
    .io_cfg_data(gibs_47_io_cfg_data),
    .io_ipinNW_0(gibs_47_io_ipinNW_0),
    .io_ipinNW_1(gibs_47_io_ipinNW_1),
    .io_opinNW_0(gibs_47_io_opinNW_0),
    .io_ipinNE_0(gibs_47_io_ipinNE_0),
    .io_ipinNE_1(gibs_47_io_ipinNE_1),
    .io_opinNE_0(gibs_47_io_opinNE_0),
    .io_ipinSE_0(gibs_47_io_ipinSE_0),
    .io_ipinSE_1(gibs_47_io_ipinSE_1),
    .io_opinSE_0(gibs_47_io_opinSE_0),
    .io_ipinSW_0(gibs_47_io_ipinSW_0),
    .io_ipinSW_1(gibs_47_io_ipinSW_1),
    .io_opinSW_0(gibs_47_io_opinSW_0),
    .io_itrackW_0(gibs_47_io_itrackW_0),
    .io_otrackW_0(gibs_47_io_otrackW_0),
    .io_itrackN_0(gibs_47_io_itrackN_0),
    .io_otrackN_0(gibs_47_io_otrackN_0),
    .io_itrackE_0(gibs_47_io_itrackE_0),
    .io_otrackE_0(gibs_47_io_otrackE_0),
    .io_itrackS_0(gibs_47_io_itrackS_0),
    .io_otrackS_0(gibs_47_io_otrackS_0)
  );
  GIB_48 gibs_48 ( // @[CGRA.scala 273:21]
    .clock(gibs_48_clock),
    .reset(gibs_48_reset),
    .io_cfg_en(gibs_48_io_cfg_en),
    .io_cfg_addr(gibs_48_io_cfg_addr),
    .io_cfg_data(gibs_48_io_cfg_data),
    .io_ipinNW_0(gibs_48_io_ipinNW_0),
    .io_ipinNW_1(gibs_48_io_ipinNW_1),
    .io_opinNW_0(gibs_48_io_opinNW_0),
    .io_ipinNE_0(gibs_48_io_ipinNE_0),
    .io_ipinNE_1(gibs_48_io_ipinNE_1),
    .io_opinNE_0(gibs_48_io_opinNE_0),
    .io_ipinSE_0(gibs_48_io_ipinSE_0),
    .io_ipinSE_1(gibs_48_io_ipinSE_1),
    .io_opinSE_0(gibs_48_io_opinSE_0),
    .io_ipinSW_0(gibs_48_io_ipinSW_0),
    .io_ipinSW_1(gibs_48_io_ipinSW_1),
    .io_opinSW_0(gibs_48_io_opinSW_0),
    .io_itrackW_0(gibs_48_io_itrackW_0),
    .io_otrackW_0(gibs_48_io_otrackW_0),
    .io_itrackN_0(gibs_48_io_itrackN_0),
    .io_otrackN_0(gibs_48_io_otrackN_0),
    .io_itrackE_0(gibs_48_io_itrackE_0),
    .io_otrackE_0(gibs_48_io_otrackE_0),
    .io_itrackS_0(gibs_48_io_itrackS_0),
    .io_otrackS_0(gibs_48_io_otrackS_0)
  );
  GIB_49 gibs_49 ( // @[CGRA.scala 273:21]
    .clock(gibs_49_clock),
    .reset(gibs_49_reset),
    .io_cfg_en(gibs_49_io_cfg_en),
    .io_cfg_addr(gibs_49_io_cfg_addr),
    .io_cfg_data(gibs_49_io_cfg_data),
    .io_ipinNW_0(gibs_49_io_ipinNW_0),
    .io_ipinNW_1(gibs_49_io_ipinNW_1),
    .io_opinNW_0(gibs_49_io_opinNW_0),
    .io_ipinNE_0(gibs_49_io_ipinNE_0),
    .io_ipinNE_1(gibs_49_io_ipinNE_1),
    .io_opinNE_0(gibs_49_io_opinNE_0),
    .io_ipinSE_0(gibs_49_io_ipinSE_0),
    .io_ipinSE_1(gibs_49_io_ipinSE_1),
    .io_opinSE_0(gibs_49_io_opinSE_0),
    .io_ipinSW_0(gibs_49_io_ipinSW_0),
    .io_ipinSW_1(gibs_49_io_ipinSW_1),
    .io_opinSW_0(gibs_49_io_opinSW_0),
    .io_itrackW_0(gibs_49_io_itrackW_0),
    .io_otrackW_0(gibs_49_io_otrackW_0),
    .io_itrackN_0(gibs_49_io_itrackN_0),
    .io_otrackN_0(gibs_49_io_otrackN_0),
    .io_itrackE_0(gibs_49_io_itrackE_0),
    .io_otrackE_0(gibs_49_io_otrackE_0),
    .io_itrackS_0(gibs_49_io_itrackS_0),
    .io_otrackS_0(gibs_49_io_otrackS_0)
  );
  GIB_50 gibs_50 ( // @[CGRA.scala 273:21]
    .clock(gibs_50_clock),
    .reset(gibs_50_reset),
    .io_cfg_en(gibs_50_io_cfg_en),
    .io_cfg_addr(gibs_50_io_cfg_addr),
    .io_cfg_data(gibs_50_io_cfg_data),
    .io_ipinNW_0(gibs_50_io_ipinNW_0),
    .io_ipinNW_1(gibs_50_io_ipinNW_1),
    .io_opinNW_0(gibs_50_io_opinNW_0),
    .io_ipinNE_0(gibs_50_io_ipinNE_0),
    .io_ipinNE_1(gibs_50_io_ipinNE_1),
    .io_opinNE_0(gibs_50_io_opinNE_0),
    .io_ipinSE_0(gibs_50_io_ipinSE_0),
    .io_ipinSE_1(gibs_50_io_ipinSE_1),
    .io_opinSE_0(gibs_50_io_opinSE_0),
    .io_ipinSW_0(gibs_50_io_ipinSW_0),
    .io_ipinSW_1(gibs_50_io_ipinSW_1),
    .io_opinSW_0(gibs_50_io_opinSW_0),
    .io_itrackW_0(gibs_50_io_itrackW_0),
    .io_otrackW_0(gibs_50_io_otrackW_0),
    .io_itrackN_0(gibs_50_io_itrackN_0),
    .io_otrackN_0(gibs_50_io_otrackN_0),
    .io_itrackE_0(gibs_50_io_itrackE_0),
    .io_otrackE_0(gibs_50_io_otrackE_0),
    .io_itrackS_0(gibs_50_io_itrackS_0),
    .io_otrackS_0(gibs_50_io_otrackS_0)
  );
  GIB_51 gibs_51 ( // @[CGRA.scala 273:21]
    .clock(gibs_51_clock),
    .reset(gibs_51_reset),
    .io_cfg_en(gibs_51_io_cfg_en),
    .io_cfg_addr(gibs_51_io_cfg_addr),
    .io_cfg_data(gibs_51_io_cfg_data),
    .io_ipinNW_0(gibs_51_io_ipinNW_0),
    .io_ipinNW_1(gibs_51_io_ipinNW_1),
    .io_opinNW_0(gibs_51_io_opinNW_0),
    .io_ipinNE_0(gibs_51_io_ipinNE_0),
    .io_ipinNE_1(gibs_51_io_ipinNE_1),
    .io_opinNE_0(gibs_51_io_opinNE_0),
    .io_ipinSE_0(gibs_51_io_ipinSE_0),
    .io_ipinSE_1(gibs_51_io_ipinSE_1),
    .io_opinSE_0(gibs_51_io_opinSE_0),
    .io_ipinSW_0(gibs_51_io_ipinSW_0),
    .io_ipinSW_1(gibs_51_io_ipinSW_1),
    .io_opinSW_0(gibs_51_io_opinSW_0),
    .io_itrackW_0(gibs_51_io_itrackW_0),
    .io_otrackW_0(gibs_51_io_otrackW_0),
    .io_itrackN_0(gibs_51_io_itrackN_0),
    .io_otrackN_0(gibs_51_io_otrackN_0),
    .io_itrackE_0(gibs_51_io_itrackE_0),
    .io_otrackE_0(gibs_51_io_otrackE_0),
    .io_itrackS_0(gibs_51_io_itrackS_0),
    .io_otrackS_0(gibs_51_io_otrackS_0)
  );
  GIB_52 gibs_52 ( // @[CGRA.scala 273:21]
    .clock(gibs_52_clock),
    .reset(gibs_52_reset),
    .io_cfg_en(gibs_52_io_cfg_en),
    .io_cfg_addr(gibs_52_io_cfg_addr),
    .io_cfg_data(gibs_52_io_cfg_data),
    .io_ipinNW_0(gibs_52_io_ipinNW_0),
    .io_ipinNW_1(gibs_52_io_ipinNW_1),
    .io_opinNW_0(gibs_52_io_opinNW_0),
    .io_ipinNE_0(gibs_52_io_ipinNE_0),
    .io_ipinNE_1(gibs_52_io_ipinNE_1),
    .io_opinNE_0(gibs_52_io_opinNE_0),
    .io_ipinSE_0(gibs_52_io_ipinSE_0),
    .io_ipinSE_1(gibs_52_io_ipinSE_1),
    .io_opinSE_0(gibs_52_io_opinSE_0),
    .io_ipinSW_0(gibs_52_io_ipinSW_0),
    .io_ipinSW_1(gibs_52_io_ipinSW_1),
    .io_opinSW_0(gibs_52_io_opinSW_0),
    .io_itrackW_0(gibs_52_io_itrackW_0),
    .io_otrackW_0(gibs_52_io_otrackW_0),
    .io_itrackN_0(gibs_52_io_itrackN_0),
    .io_otrackN_0(gibs_52_io_otrackN_0),
    .io_itrackE_0(gibs_52_io_itrackE_0),
    .io_otrackE_0(gibs_52_io_otrackE_0),
    .io_itrackS_0(gibs_52_io_itrackS_0),
    .io_otrackS_0(gibs_52_io_otrackS_0)
  );
  GIB_53 gibs_53 ( // @[CGRA.scala 273:21]
    .clock(gibs_53_clock),
    .reset(gibs_53_reset),
    .io_cfg_en(gibs_53_io_cfg_en),
    .io_cfg_addr(gibs_53_io_cfg_addr),
    .io_cfg_data(gibs_53_io_cfg_data),
    .io_ipinNW_0(gibs_53_io_ipinNW_0),
    .io_ipinNW_1(gibs_53_io_ipinNW_1),
    .io_opinNW_0(gibs_53_io_opinNW_0),
    .io_ipinSW_0(gibs_53_io_ipinSW_0),
    .io_ipinSW_1(gibs_53_io_ipinSW_1),
    .io_opinSW_0(gibs_53_io_opinSW_0),
    .io_itrackW_0(gibs_53_io_itrackW_0),
    .io_otrackW_0(gibs_53_io_otrackW_0),
    .io_itrackN_0(gibs_53_io_itrackN_0),
    .io_otrackN_0(gibs_53_io_otrackN_0),
    .io_itrackS_0(gibs_53_io_itrackS_0),
    .io_otrackS_0(gibs_53_io_otrackS_0)
  );
  GIB_54 gibs_54 ( // @[CGRA.scala 273:21]
    .clock(gibs_54_clock),
    .reset(gibs_54_reset),
    .io_cfg_en(gibs_54_io_cfg_en),
    .io_cfg_addr(gibs_54_io_cfg_addr),
    .io_cfg_data(gibs_54_io_cfg_data),
    .io_ipinNE_0(gibs_54_io_ipinNE_0),
    .io_ipinNE_1(gibs_54_io_ipinNE_1),
    .io_opinNE_0(gibs_54_io_opinNE_0),
    .io_ipinSE_0(gibs_54_io_ipinSE_0),
    .io_ipinSE_1(gibs_54_io_ipinSE_1),
    .io_opinSE_0(gibs_54_io_opinSE_0),
    .io_itrackN_0(gibs_54_io_itrackN_0),
    .io_otrackN_0(gibs_54_io_otrackN_0),
    .io_itrackE_0(gibs_54_io_itrackE_0),
    .io_otrackE_0(gibs_54_io_otrackE_0),
    .io_itrackS_0(gibs_54_io_itrackS_0),
    .io_otrackS_0(gibs_54_io_otrackS_0)
  );
  GIB_55 gibs_55 ( // @[CGRA.scala 273:21]
    .clock(gibs_55_clock),
    .reset(gibs_55_reset),
    .io_cfg_en(gibs_55_io_cfg_en),
    .io_cfg_addr(gibs_55_io_cfg_addr),
    .io_cfg_data(gibs_55_io_cfg_data),
    .io_ipinNW_0(gibs_55_io_ipinNW_0),
    .io_ipinNW_1(gibs_55_io_ipinNW_1),
    .io_opinNW_0(gibs_55_io_opinNW_0),
    .io_ipinNE_0(gibs_55_io_ipinNE_0),
    .io_ipinNE_1(gibs_55_io_ipinNE_1),
    .io_opinNE_0(gibs_55_io_opinNE_0),
    .io_ipinSE_0(gibs_55_io_ipinSE_0),
    .io_ipinSE_1(gibs_55_io_ipinSE_1),
    .io_opinSE_0(gibs_55_io_opinSE_0),
    .io_ipinSW_0(gibs_55_io_ipinSW_0),
    .io_ipinSW_1(gibs_55_io_ipinSW_1),
    .io_opinSW_0(gibs_55_io_opinSW_0),
    .io_itrackW_0(gibs_55_io_itrackW_0),
    .io_otrackW_0(gibs_55_io_otrackW_0),
    .io_itrackN_0(gibs_55_io_itrackN_0),
    .io_otrackN_0(gibs_55_io_otrackN_0),
    .io_itrackE_0(gibs_55_io_itrackE_0),
    .io_otrackE_0(gibs_55_io_otrackE_0),
    .io_itrackS_0(gibs_55_io_itrackS_0),
    .io_otrackS_0(gibs_55_io_otrackS_0)
  );
  GIB_56 gibs_56 ( // @[CGRA.scala 273:21]
    .clock(gibs_56_clock),
    .reset(gibs_56_reset),
    .io_cfg_en(gibs_56_io_cfg_en),
    .io_cfg_addr(gibs_56_io_cfg_addr),
    .io_cfg_data(gibs_56_io_cfg_data),
    .io_ipinNW_0(gibs_56_io_ipinNW_0),
    .io_ipinNW_1(gibs_56_io_ipinNW_1),
    .io_opinNW_0(gibs_56_io_opinNW_0),
    .io_ipinNE_0(gibs_56_io_ipinNE_0),
    .io_ipinNE_1(gibs_56_io_ipinNE_1),
    .io_opinNE_0(gibs_56_io_opinNE_0),
    .io_ipinSE_0(gibs_56_io_ipinSE_0),
    .io_ipinSE_1(gibs_56_io_ipinSE_1),
    .io_opinSE_0(gibs_56_io_opinSE_0),
    .io_ipinSW_0(gibs_56_io_ipinSW_0),
    .io_ipinSW_1(gibs_56_io_ipinSW_1),
    .io_opinSW_0(gibs_56_io_opinSW_0),
    .io_itrackW_0(gibs_56_io_itrackW_0),
    .io_otrackW_0(gibs_56_io_otrackW_0),
    .io_itrackN_0(gibs_56_io_itrackN_0),
    .io_otrackN_0(gibs_56_io_otrackN_0),
    .io_itrackE_0(gibs_56_io_itrackE_0),
    .io_otrackE_0(gibs_56_io_otrackE_0),
    .io_itrackS_0(gibs_56_io_itrackS_0),
    .io_otrackS_0(gibs_56_io_otrackS_0)
  );
  GIB_57 gibs_57 ( // @[CGRA.scala 273:21]
    .clock(gibs_57_clock),
    .reset(gibs_57_reset),
    .io_cfg_en(gibs_57_io_cfg_en),
    .io_cfg_addr(gibs_57_io_cfg_addr),
    .io_cfg_data(gibs_57_io_cfg_data),
    .io_ipinNW_0(gibs_57_io_ipinNW_0),
    .io_ipinNW_1(gibs_57_io_ipinNW_1),
    .io_opinNW_0(gibs_57_io_opinNW_0),
    .io_ipinNE_0(gibs_57_io_ipinNE_0),
    .io_ipinNE_1(gibs_57_io_ipinNE_1),
    .io_opinNE_0(gibs_57_io_opinNE_0),
    .io_ipinSE_0(gibs_57_io_ipinSE_0),
    .io_ipinSE_1(gibs_57_io_ipinSE_1),
    .io_opinSE_0(gibs_57_io_opinSE_0),
    .io_ipinSW_0(gibs_57_io_ipinSW_0),
    .io_ipinSW_1(gibs_57_io_ipinSW_1),
    .io_opinSW_0(gibs_57_io_opinSW_0),
    .io_itrackW_0(gibs_57_io_itrackW_0),
    .io_otrackW_0(gibs_57_io_otrackW_0),
    .io_itrackN_0(gibs_57_io_itrackN_0),
    .io_otrackN_0(gibs_57_io_otrackN_0),
    .io_itrackE_0(gibs_57_io_itrackE_0),
    .io_otrackE_0(gibs_57_io_otrackE_0),
    .io_itrackS_0(gibs_57_io_itrackS_0),
    .io_otrackS_0(gibs_57_io_otrackS_0)
  );
  GIB_58 gibs_58 ( // @[CGRA.scala 273:21]
    .clock(gibs_58_clock),
    .reset(gibs_58_reset),
    .io_cfg_en(gibs_58_io_cfg_en),
    .io_cfg_addr(gibs_58_io_cfg_addr),
    .io_cfg_data(gibs_58_io_cfg_data),
    .io_ipinNW_0(gibs_58_io_ipinNW_0),
    .io_ipinNW_1(gibs_58_io_ipinNW_1),
    .io_opinNW_0(gibs_58_io_opinNW_0),
    .io_ipinNE_0(gibs_58_io_ipinNE_0),
    .io_ipinNE_1(gibs_58_io_ipinNE_1),
    .io_opinNE_0(gibs_58_io_opinNE_0),
    .io_ipinSE_0(gibs_58_io_ipinSE_0),
    .io_ipinSE_1(gibs_58_io_ipinSE_1),
    .io_opinSE_0(gibs_58_io_opinSE_0),
    .io_ipinSW_0(gibs_58_io_ipinSW_0),
    .io_ipinSW_1(gibs_58_io_ipinSW_1),
    .io_opinSW_0(gibs_58_io_opinSW_0),
    .io_itrackW_0(gibs_58_io_itrackW_0),
    .io_otrackW_0(gibs_58_io_otrackW_0),
    .io_itrackN_0(gibs_58_io_itrackN_0),
    .io_otrackN_0(gibs_58_io_otrackN_0),
    .io_itrackE_0(gibs_58_io_itrackE_0),
    .io_otrackE_0(gibs_58_io_otrackE_0),
    .io_itrackS_0(gibs_58_io_itrackS_0),
    .io_otrackS_0(gibs_58_io_otrackS_0)
  );
  GIB_59 gibs_59 ( // @[CGRA.scala 273:21]
    .clock(gibs_59_clock),
    .reset(gibs_59_reset),
    .io_cfg_en(gibs_59_io_cfg_en),
    .io_cfg_addr(gibs_59_io_cfg_addr),
    .io_cfg_data(gibs_59_io_cfg_data),
    .io_ipinNW_0(gibs_59_io_ipinNW_0),
    .io_ipinNW_1(gibs_59_io_ipinNW_1),
    .io_opinNW_0(gibs_59_io_opinNW_0),
    .io_ipinNE_0(gibs_59_io_ipinNE_0),
    .io_ipinNE_1(gibs_59_io_ipinNE_1),
    .io_opinNE_0(gibs_59_io_opinNE_0),
    .io_ipinSE_0(gibs_59_io_ipinSE_0),
    .io_ipinSE_1(gibs_59_io_ipinSE_1),
    .io_opinSE_0(gibs_59_io_opinSE_0),
    .io_ipinSW_0(gibs_59_io_ipinSW_0),
    .io_ipinSW_1(gibs_59_io_ipinSW_1),
    .io_opinSW_0(gibs_59_io_opinSW_0),
    .io_itrackW_0(gibs_59_io_itrackW_0),
    .io_otrackW_0(gibs_59_io_otrackW_0),
    .io_itrackN_0(gibs_59_io_itrackN_0),
    .io_otrackN_0(gibs_59_io_otrackN_0),
    .io_itrackE_0(gibs_59_io_itrackE_0),
    .io_otrackE_0(gibs_59_io_otrackE_0),
    .io_itrackS_0(gibs_59_io_itrackS_0),
    .io_otrackS_0(gibs_59_io_otrackS_0)
  );
  GIB_60 gibs_60 ( // @[CGRA.scala 273:21]
    .clock(gibs_60_clock),
    .reset(gibs_60_reset),
    .io_cfg_en(gibs_60_io_cfg_en),
    .io_cfg_addr(gibs_60_io_cfg_addr),
    .io_cfg_data(gibs_60_io_cfg_data),
    .io_ipinNW_0(gibs_60_io_ipinNW_0),
    .io_ipinNW_1(gibs_60_io_ipinNW_1),
    .io_opinNW_0(gibs_60_io_opinNW_0),
    .io_ipinNE_0(gibs_60_io_ipinNE_0),
    .io_ipinNE_1(gibs_60_io_ipinNE_1),
    .io_opinNE_0(gibs_60_io_opinNE_0),
    .io_ipinSE_0(gibs_60_io_ipinSE_0),
    .io_ipinSE_1(gibs_60_io_ipinSE_1),
    .io_opinSE_0(gibs_60_io_opinSE_0),
    .io_ipinSW_0(gibs_60_io_ipinSW_0),
    .io_ipinSW_1(gibs_60_io_ipinSW_1),
    .io_opinSW_0(gibs_60_io_opinSW_0),
    .io_itrackW_0(gibs_60_io_itrackW_0),
    .io_otrackW_0(gibs_60_io_otrackW_0),
    .io_itrackN_0(gibs_60_io_itrackN_0),
    .io_otrackN_0(gibs_60_io_otrackN_0),
    .io_itrackE_0(gibs_60_io_itrackE_0),
    .io_otrackE_0(gibs_60_io_otrackE_0),
    .io_itrackS_0(gibs_60_io_itrackS_0),
    .io_otrackS_0(gibs_60_io_otrackS_0)
  );
  GIB_61 gibs_61 ( // @[CGRA.scala 273:21]
    .clock(gibs_61_clock),
    .reset(gibs_61_reset),
    .io_cfg_en(gibs_61_io_cfg_en),
    .io_cfg_addr(gibs_61_io_cfg_addr),
    .io_cfg_data(gibs_61_io_cfg_data),
    .io_ipinNW_0(gibs_61_io_ipinNW_0),
    .io_ipinNW_1(gibs_61_io_ipinNW_1),
    .io_opinNW_0(gibs_61_io_opinNW_0),
    .io_ipinNE_0(gibs_61_io_ipinNE_0),
    .io_ipinNE_1(gibs_61_io_ipinNE_1),
    .io_opinNE_0(gibs_61_io_opinNE_0),
    .io_ipinSE_0(gibs_61_io_ipinSE_0),
    .io_ipinSE_1(gibs_61_io_ipinSE_1),
    .io_opinSE_0(gibs_61_io_opinSE_0),
    .io_ipinSW_0(gibs_61_io_ipinSW_0),
    .io_ipinSW_1(gibs_61_io_ipinSW_1),
    .io_opinSW_0(gibs_61_io_opinSW_0),
    .io_itrackW_0(gibs_61_io_itrackW_0),
    .io_otrackW_0(gibs_61_io_otrackW_0),
    .io_itrackN_0(gibs_61_io_itrackN_0),
    .io_otrackN_0(gibs_61_io_otrackN_0),
    .io_itrackE_0(gibs_61_io_itrackE_0),
    .io_otrackE_0(gibs_61_io_otrackE_0),
    .io_itrackS_0(gibs_61_io_itrackS_0),
    .io_otrackS_0(gibs_61_io_otrackS_0)
  );
  GIB_62 gibs_62 ( // @[CGRA.scala 273:21]
    .clock(gibs_62_clock),
    .reset(gibs_62_reset),
    .io_cfg_en(gibs_62_io_cfg_en),
    .io_cfg_addr(gibs_62_io_cfg_addr),
    .io_cfg_data(gibs_62_io_cfg_data),
    .io_ipinNW_0(gibs_62_io_ipinNW_0),
    .io_ipinNW_1(gibs_62_io_ipinNW_1),
    .io_opinNW_0(gibs_62_io_opinNW_0),
    .io_ipinSW_0(gibs_62_io_ipinSW_0),
    .io_ipinSW_1(gibs_62_io_ipinSW_1),
    .io_opinSW_0(gibs_62_io_opinSW_0),
    .io_itrackW_0(gibs_62_io_itrackW_0),
    .io_otrackW_0(gibs_62_io_otrackW_0),
    .io_itrackN_0(gibs_62_io_itrackN_0),
    .io_otrackN_0(gibs_62_io_otrackN_0),
    .io_itrackS_0(gibs_62_io_itrackS_0),
    .io_otrackS_0(gibs_62_io_otrackS_0)
  );
  GIB_63 gibs_63 ( // @[CGRA.scala 273:21]
    .clock(gibs_63_clock),
    .reset(gibs_63_reset),
    .io_cfg_en(gibs_63_io_cfg_en),
    .io_cfg_addr(gibs_63_io_cfg_addr),
    .io_cfg_data(gibs_63_io_cfg_data),
    .io_ipinNE_0(gibs_63_io_ipinNE_0),
    .io_ipinNE_1(gibs_63_io_ipinNE_1),
    .io_opinNE_0(gibs_63_io_opinNE_0),
    .io_ipinSE_0(gibs_63_io_ipinSE_0),
    .io_ipinSE_1(gibs_63_io_ipinSE_1),
    .io_opinSE_0(gibs_63_io_opinSE_0),
    .io_itrackN_0(gibs_63_io_itrackN_0),
    .io_otrackN_0(gibs_63_io_otrackN_0),
    .io_itrackE_0(gibs_63_io_itrackE_0),
    .io_otrackE_0(gibs_63_io_otrackE_0),
    .io_itrackS_0(gibs_63_io_itrackS_0),
    .io_otrackS_0(gibs_63_io_otrackS_0)
  );
  GIB_64 gibs_64 ( // @[CGRA.scala 273:21]
    .clock(gibs_64_clock),
    .reset(gibs_64_reset),
    .io_cfg_en(gibs_64_io_cfg_en),
    .io_cfg_addr(gibs_64_io_cfg_addr),
    .io_cfg_data(gibs_64_io_cfg_data),
    .io_ipinNW_0(gibs_64_io_ipinNW_0),
    .io_ipinNW_1(gibs_64_io_ipinNW_1),
    .io_opinNW_0(gibs_64_io_opinNW_0),
    .io_ipinNE_0(gibs_64_io_ipinNE_0),
    .io_ipinNE_1(gibs_64_io_ipinNE_1),
    .io_opinNE_0(gibs_64_io_opinNE_0),
    .io_ipinSE_0(gibs_64_io_ipinSE_0),
    .io_ipinSE_1(gibs_64_io_ipinSE_1),
    .io_opinSE_0(gibs_64_io_opinSE_0),
    .io_ipinSW_0(gibs_64_io_ipinSW_0),
    .io_ipinSW_1(gibs_64_io_ipinSW_1),
    .io_opinSW_0(gibs_64_io_opinSW_0),
    .io_itrackW_0(gibs_64_io_itrackW_0),
    .io_otrackW_0(gibs_64_io_otrackW_0),
    .io_itrackN_0(gibs_64_io_itrackN_0),
    .io_otrackN_0(gibs_64_io_otrackN_0),
    .io_itrackE_0(gibs_64_io_itrackE_0),
    .io_otrackE_0(gibs_64_io_otrackE_0),
    .io_itrackS_0(gibs_64_io_itrackS_0),
    .io_otrackS_0(gibs_64_io_otrackS_0)
  );
  GIB_65 gibs_65 ( // @[CGRA.scala 273:21]
    .clock(gibs_65_clock),
    .reset(gibs_65_reset),
    .io_cfg_en(gibs_65_io_cfg_en),
    .io_cfg_addr(gibs_65_io_cfg_addr),
    .io_cfg_data(gibs_65_io_cfg_data),
    .io_ipinNW_0(gibs_65_io_ipinNW_0),
    .io_ipinNW_1(gibs_65_io_ipinNW_1),
    .io_opinNW_0(gibs_65_io_opinNW_0),
    .io_ipinNE_0(gibs_65_io_ipinNE_0),
    .io_ipinNE_1(gibs_65_io_ipinNE_1),
    .io_opinNE_0(gibs_65_io_opinNE_0),
    .io_ipinSE_0(gibs_65_io_ipinSE_0),
    .io_ipinSE_1(gibs_65_io_ipinSE_1),
    .io_opinSE_0(gibs_65_io_opinSE_0),
    .io_ipinSW_0(gibs_65_io_ipinSW_0),
    .io_ipinSW_1(gibs_65_io_ipinSW_1),
    .io_opinSW_0(gibs_65_io_opinSW_0),
    .io_itrackW_0(gibs_65_io_itrackW_0),
    .io_otrackW_0(gibs_65_io_otrackW_0),
    .io_itrackN_0(gibs_65_io_itrackN_0),
    .io_otrackN_0(gibs_65_io_otrackN_0),
    .io_itrackE_0(gibs_65_io_itrackE_0),
    .io_otrackE_0(gibs_65_io_otrackE_0),
    .io_itrackS_0(gibs_65_io_itrackS_0),
    .io_otrackS_0(gibs_65_io_otrackS_0)
  );
  GIB_66 gibs_66 ( // @[CGRA.scala 273:21]
    .clock(gibs_66_clock),
    .reset(gibs_66_reset),
    .io_cfg_en(gibs_66_io_cfg_en),
    .io_cfg_addr(gibs_66_io_cfg_addr),
    .io_cfg_data(gibs_66_io_cfg_data),
    .io_ipinNW_0(gibs_66_io_ipinNW_0),
    .io_ipinNW_1(gibs_66_io_ipinNW_1),
    .io_opinNW_0(gibs_66_io_opinNW_0),
    .io_ipinNE_0(gibs_66_io_ipinNE_0),
    .io_ipinNE_1(gibs_66_io_ipinNE_1),
    .io_opinNE_0(gibs_66_io_opinNE_0),
    .io_ipinSE_0(gibs_66_io_ipinSE_0),
    .io_ipinSE_1(gibs_66_io_ipinSE_1),
    .io_opinSE_0(gibs_66_io_opinSE_0),
    .io_ipinSW_0(gibs_66_io_ipinSW_0),
    .io_ipinSW_1(gibs_66_io_ipinSW_1),
    .io_opinSW_0(gibs_66_io_opinSW_0),
    .io_itrackW_0(gibs_66_io_itrackW_0),
    .io_otrackW_0(gibs_66_io_otrackW_0),
    .io_itrackN_0(gibs_66_io_itrackN_0),
    .io_otrackN_0(gibs_66_io_otrackN_0),
    .io_itrackE_0(gibs_66_io_itrackE_0),
    .io_otrackE_0(gibs_66_io_otrackE_0),
    .io_itrackS_0(gibs_66_io_itrackS_0),
    .io_otrackS_0(gibs_66_io_otrackS_0)
  );
  GIB_67 gibs_67 ( // @[CGRA.scala 273:21]
    .clock(gibs_67_clock),
    .reset(gibs_67_reset),
    .io_cfg_en(gibs_67_io_cfg_en),
    .io_cfg_addr(gibs_67_io_cfg_addr),
    .io_cfg_data(gibs_67_io_cfg_data),
    .io_ipinNW_0(gibs_67_io_ipinNW_0),
    .io_ipinNW_1(gibs_67_io_ipinNW_1),
    .io_opinNW_0(gibs_67_io_opinNW_0),
    .io_ipinNE_0(gibs_67_io_ipinNE_0),
    .io_ipinNE_1(gibs_67_io_ipinNE_1),
    .io_opinNE_0(gibs_67_io_opinNE_0),
    .io_ipinSE_0(gibs_67_io_ipinSE_0),
    .io_ipinSE_1(gibs_67_io_ipinSE_1),
    .io_opinSE_0(gibs_67_io_opinSE_0),
    .io_ipinSW_0(gibs_67_io_ipinSW_0),
    .io_ipinSW_1(gibs_67_io_ipinSW_1),
    .io_opinSW_0(gibs_67_io_opinSW_0),
    .io_itrackW_0(gibs_67_io_itrackW_0),
    .io_otrackW_0(gibs_67_io_otrackW_0),
    .io_itrackN_0(gibs_67_io_itrackN_0),
    .io_otrackN_0(gibs_67_io_otrackN_0),
    .io_itrackE_0(gibs_67_io_itrackE_0),
    .io_otrackE_0(gibs_67_io_otrackE_0),
    .io_itrackS_0(gibs_67_io_itrackS_0),
    .io_otrackS_0(gibs_67_io_otrackS_0)
  );
  GIB_68 gibs_68 ( // @[CGRA.scala 273:21]
    .clock(gibs_68_clock),
    .reset(gibs_68_reset),
    .io_cfg_en(gibs_68_io_cfg_en),
    .io_cfg_addr(gibs_68_io_cfg_addr),
    .io_cfg_data(gibs_68_io_cfg_data),
    .io_ipinNW_0(gibs_68_io_ipinNW_0),
    .io_ipinNW_1(gibs_68_io_ipinNW_1),
    .io_opinNW_0(gibs_68_io_opinNW_0),
    .io_ipinNE_0(gibs_68_io_ipinNE_0),
    .io_ipinNE_1(gibs_68_io_ipinNE_1),
    .io_opinNE_0(gibs_68_io_opinNE_0),
    .io_ipinSE_0(gibs_68_io_ipinSE_0),
    .io_ipinSE_1(gibs_68_io_ipinSE_1),
    .io_opinSE_0(gibs_68_io_opinSE_0),
    .io_ipinSW_0(gibs_68_io_ipinSW_0),
    .io_ipinSW_1(gibs_68_io_ipinSW_1),
    .io_opinSW_0(gibs_68_io_opinSW_0),
    .io_itrackW_0(gibs_68_io_itrackW_0),
    .io_otrackW_0(gibs_68_io_otrackW_0),
    .io_itrackN_0(gibs_68_io_itrackN_0),
    .io_otrackN_0(gibs_68_io_otrackN_0),
    .io_itrackE_0(gibs_68_io_itrackE_0),
    .io_otrackE_0(gibs_68_io_otrackE_0),
    .io_itrackS_0(gibs_68_io_itrackS_0),
    .io_otrackS_0(gibs_68_io_otrackS_0)
  );
  GIB_69 gibs_69 ( // @[CGRA.scala 273:21]
    .clock(gibs_69_clock),
    .reset(gibs_69_reset),
    .io_cfg_en(gibs_69_io_cfg_en),
    .io_cfg_addr(gibs_69_io_cfg_addr),
    .io_cfg_data(gibs_69_io_cfg_data),
    .io_ipinNW_0(gibs_69_io_ipinNW_0),
    .io_ipinNW_1(gibs_69_io_ipinNW_1),
    .io_opinNW_0(gibs_69_io_opinNW_0),
    .io_ipinNE_0(gibs_69_io_ipinNE_0),
    .io_ipinNE_1(gibs_69_io_ipinNE_1),
    .io_opinNE_0(gibs_69_io_opinNE_0),
    .io_ipinSE_0(gibs_69_io_ipinSE_0),
    .io_ipinSE_1(gibs_69_io_ipinSE_1),
    .io_opinSE_0(gibs_69_io_opinSE_0),
    .io_ipinSW_0(gibs_69_io_ipinSW_0),
    .io_ipinSW_1(gibs_69_io_ipinSW_1),
    .io_opinSW_0(gibs_69_io_opinSW_0),
    .io_itrackW_0(gibs_69_io_itrackW_0),
    .io_otrackW_0(gibs_69_io_otrackW_0),
    .io_itrackN_0(gibs_69_io_itrackN_0),
    .io_otrackN_0(gibs_69_io_otrackN_0),
    .io_itrackE_0(gibs_69_io_itrackE_0),
    .io_otrackE_0(gibs_69_io_otrackE_0),
    .io_itrackS_0(gibs_69_io_itrackS_0),
    .io_otrackS_0(gibs_69_io_otrackS_0)
  );
  GIB_70 gibs_70 ( // @[CGRA.scala 273:21]
    .clock(gibs_70_clock),
    .reset(gibs_70_reset),
    .io_cfg_en(gibs_70_io_cfg_en),
    .io_cfg_addr(gibs_70_io_cfg_addr),
    .io_cfg_data(gibs_70_io_cfg_data),
    .io_ipinNW_0(gibs_70_io_ipinNW_0),
    .io_ipinNW_1(gibs_70_io_ipinNW_1),
    .io_opinNW_0(gibs_70_io_opinNW_0),
    .io_ipinNE_0(gibs_70_io_ipinNE_0),
    .io_ipinNE_1(gibs_70_io_ipinNE_1),
    .io_opinNE_0(gibs_70_io_opinNE_0),
    .io_ipinSE_0(gibs_70_io_ipinSE_0),
    .io_ipinSE_1(gibs_70_io_ipinSE_1),
    .io_opinSE_0(gibs_70_io_opinSE_0),
    .io_ipinSW_0(gibs_70_io_ipinSW_0),
    .io_ipinSW_1(gibs_70_io_ipinSW_1),
    .io_opinSW_0(gibs_70_io_opinSW_0),
    .io_itrackW_0(gibs_70_io_itrackW_0),
    .io_otrackW_0(gibs_70_io_otrackW_0),
    .io_itrackN_0(gibs_70_io_itrackN_0),
    .io_otrackN_0(gibs_70_io_otrackN_0),
    .io_itrackE_0(gibs_70_io_itrackE_0),
    .io_otrackE_0(gibs_70_io_otrackE_0),
    .io_itrackS_0(gibs_70_io_itrackS_0),
    .io_otrackS_0(gibs_70_io_otrackS_0)
  );
  GIB_71 gibs_71 ( // @[CGRA.scala 273:21]
    .clock(gibs_71_clock),
    .reset(gibs_71_reset),
    .io_cfg_en(gibs_71_io_cfg_en),
    .io_cfg_addr(gibs_71_io_cfg_addr),
    .io_cfg_data(gibs_71_io_cfg_data),
    .io_ipinNW_0(gibs_71_io_ipinNW_0),
    .io_ipinNW_1(gibs_71_io_ipinNW_1),
    .io_opinNW_0(gibs_71_io_opinNW_0),
    .io_ipinSW_0(gibs_71_io_ipinSW_0),
    .io_ipinSW_1(gibs_71_io_ipinSW_1),
    .io_opinSW_0(gibs_71_io_opinSW_0),
    .io_itrackW_0(gibs_71_io_itrackW_0),
    .io_otrackW_0(gibs_71_io_otrackW_0),
    .io_itrackN_0(gibs_71_io_itrackN_0),
    .io_otrackN_0(gibs_71_io_otrackN_0),
    .io_itrackS_0(gibs_71_io_itrackS_0),
    .io_otrackS_0(gibs_71_io_otrackS_0)
  );
  GIB_72 gibs_72 ( // @[CGRA.scala 273:21]
    .clock(gibs_72_clock),
    .reset(gibs_72_reset),
    .io_cfg_en(gibs_72_io_cfg_en),
    .io_cfg_addr(gibs_72_io_cfg_addr),
    .io_cfg_data(gibs_72_io_cfg_data),
    .io_ipinNE_0(gibs_72_io_ipinNE_0),
    .io_ipinNE_1(gibs_72_io_ipinNE_1),
    .io_opinNE_0(gibs_72_io_opinNE_0),
    .io_ipinSE_0(gibs_72_io_ipinSE_0),
    .io_opinSE_0(gibs_72_io_opinSE_0),
    .io_itrackN_0(gibs_72_io_itrackN_0),
    .io_otrackN_0(gibs_72_io_otrackN_0),
    .io_itrackE_0(gibs_72_io_itrackE_0),
    .io_otrackE_0(gibs_72_io_otrackE_0)
  );
  GIB_73 gibs_73 ( // @[CGRA.scala 273:21]
    .clock(gibs_73_clock),
    .reset(gibs_73_reset),
    .io_cfg_en(gibs_73_io_cfg_en),
    .io_cfg_addr(gibs_73_io_cfg_addr),
    .io_cfg_data(gibs_73_io_cfg_data),
    .io_ipinNW_0(gibs_73_io_ipinNW_0),
    .io_ipinNW_1(gibs_73_io_ipinNW_1),
    .io_opinNW_0(gibs_73_io_opinNW_0),
    .io_ipinNE_0(gibs_73_io_ipinNE_0),
    .io_ipinNE_1(gibs_73_io_ipinNE_1),
    .io_opinNE_0(gibs_73_io_opinNE_0),
    .io_ipinSE_0(gibs_73_io_ipinSE_0),
    .io_opinSE_0(gibs_73_io_opinSE_0),
    .io_ipinSW_0(gibs_73_io_ipinSW_0),
    .io_opinSW_0(gibs_73_io_opinSW_0),
    .io_itrackW_0(gibs_73_io_itrackW_0),
    .io_otrackW_0(gibs_73_io_otrackW_0),
    .io_itrackN_0(gibs_73_io_itrackN_0),
    .io_otrackN_0(gibs_73_io_otrackN_0),
    .io_itrackE_0(gibs_73_io_itrackE_0),
    .io_otrackE_0(gibs_73_io_otrackE_0)
  );
  GIB_74 gibs_74 ( // @[CGRA.scala 273:21]
    .clock(gibs_74_clock),
    .reset(gibs_74_reset),
    .io_cfg_en(gibs_74_io_cfg_en),
    .io_cfg_addr(gibs_74_io_cfg_addr),
    .io_cfg_data(gibs_74_io_cfg_data),
    .io_ipinNW_0(gibs_74_io_ipinNW_0),
    .io_ipinNW_1(gibs_74_io_ipinNW_1),
    .io_opinNW_0(gibs_74_io_opinNW_0),
    .io_ipinNE_0(gibs_74_io_ipinNE_0),
    .io_ipinNE_1(gibs_74_io_ipinNE_1),
    .io_opinNE_0(gibs_74_io_opinNE_0),
    .io_ipinSE_0(gibs_74_io_ipinSE_0),
    .io_opinSE_0(gibs_74_io_opinSE_0),
    .io_ipinSW_0(gibs_74_io_ipinSW_0),
    .io_opinSW_0(gibs_74_io_opinSW_0),
    .io_itrackW_0(gibs_74_io_itrackW_0),
    .io_otrackW_0(gibs_74_io_otrackW_0),
    .io_itrackN_0(gibs_74_io_itrackN_0),
    .io_otrackN_0(gibs_74_io_otrackN_0),
    .io_itrackE_0(gibs_74_io_itrackE_0),
    .io_otrackE_0(gibs_74_io_otrackE_0)
  );
  GIB_75 gibs_75 ( // @[CGRA.scala 273:21]
    .clock(gibs_75_clock),
    .reset(gibs_75_reset),
    .io_cfg_en(gibs_75_io_cfg_en),
    .io_cfg_addr(gibs_75_io_cfg_addr),
    .io_cfg_data(gibs_75_io_cfg_data),
    .io_ipinNW_0(gibs_75_io_ipinNW_0),
    .io_ipinNW_1(gibs_75_io_ipinNW_1),
    .io_opinNW_0(gibs_75_io_opinNW_0),
    .io_ipinNE_0(gibs_75_io_ipinNE_0),
    .io_ipinNE_1(gibs_75_io_ipinNE_1),
    .io_opinNE_0(gibs_75_io_opinNE_0),
    .io_ipinSE_0(gibs_75_io_ipinSE_0),
    .io_opinSE_0(gibs_75_io_opinSE_0),
    .io_ipinSW_0(gibs_75_io_ipinSW_0),
    .io_opinSW_0(gibs_75_io_opinSW_0),
    .io_itrackW_0(gibs_75_io_itrackW_0),
    .io_otrackW_0(gibs_75_io_otrackW_0),
    .io_itrackN_0(gibs_75_io_itrackN_0),
    .io_otrackN_0(gibs_75_io_otrackN_0),
    .io_itrackE_0(gibs_75_io_itrackE_0),
    .io_otrackE_0(gibs_75_io_otrackE_0)
  );
  GIB_76 gibs_76 ( // @[CGRA.scala 273:21]
    .clock(gibs_76_clock),
    .reset(gibs_76_reset),
    .io_cfg_en(gibs_76_io_cfg_en),
    .io_cfg_addr(gibs_76_io_cfg_addr),
    .io_cfg_data(gibs_76_io_cfg_data),
    .io_ipinNW_0(gibs_76_io_ipinNW_0),
    .io_ipinNW_1(gibs_76_io_ipinNW_1),
    .io_opinNW_0(gibs_76_io_opinNW_0),
    .io_ipinNE_0(gibs_76_io_ipinNE_0),
    .io_ipinNE_1(gibs_76_io_ipinNE_1),
    .io_opinNE_0(gibs_76_io_opinNE_0),
    .io_ipinSE_0(gibs_76_io_ipinSE_0),
    .io_opinSE_0(gibs_76_io_opinSE_0),
    .io_ipinSW_0(gibs_76_io_ipinSW_0),
    .io_opinSW_0(gibs_76_io_opinSW_0),
    .io_itrackW_0(gibs_76_io_itrackW_0),
    .io_otrackW_0(gibs_76_io_otrackW_0),
    .io_itrackN_0(gibs_76_io_itrackN_0),
    .io_otrackN_0(gibs_76_io_otrackN_0),
    .io_itrackE_0(gibs_76_io_itrackE_0),
    .io_otrackE_0(gibs_76_io_otrackE_0)
  );
  GIB_77 gibs_77 ( // @[CGRA.scala 273:21]
    .clock(gibs_77_clock),
    .reset(gibs_77_reset),
    .io_cfg_en(gibs_77_io_cfg_en),
    .io_cfg_addr(gibs_77_io_cfg_addr),
    .io_cfg_data(gibs_77_io_cfg_data),
    .io_ipinNW_0(gibs_77_io_ipinNW_0),
    .io_ipinNW_1(gibs_77_io_ipinNW_1),
    .io_opinNW_0(gibs_77_io_opinNW_0),
    .io_ipinNE_0(gibs_77_io_ipinNE_0),
    .io_ipinNE_1(gibs_77_io_ipinNE_1),
    .io_opinNE_0(gibs_77_io_opinNE_0),
    .io_ipinSE_0(gibs_77_io_ipinSE_0),
    .io_opinSE_0(gibs_77_io_opinSE_0),
    .io_ipinSW_0(gibs_77_io_ipinSW_0),
    .io_opinSW_0(gibs_77_io_opinSW_0),
    .io_itrackW_0(gibs_77_io_itrackW_0),
    .io_otrackW_0(gibs_77_io_otrackW_0),
    .io_itrackN_0(gibs_77_io_itrackN_0),
    .io_otrackN_0(gibs_77_io_otrackN_0),
    .io_itrackE_0(gibs_77_io_itrackE_0),
    .io_otrackE_0(gibs_77_io_otrackE_0)
  );
  GIB_78 gibs_78 ( // @[CGRA.scala 273:21]
    .clock(gibs_78_clock),
    .reset(gibs_78_reset),
    .io_cfg_en(gibs_78_io_cfg_en),
    .io_cfg_addr(gibs_78_io_cfg_addr),
    .io_cfg_data(gibs_78_io_cfg_data),
    .io_ipinNW_0(gibs_78_io_ipinNW_0),
    .io_ipinNW_1(gibs_78_io_ipinNW_1),
    .io_opinNW_0(gibs_78_io_opinNW_0),
    .io_ipinNE_0(gibs_78_io_ipinNE_0),
    .io_ipinNE_1(gibs_78_io_ipinNE_1),
    .io_opinNE_0(gibs_78_io_opinNE_0),
    .io_ipinSE_0(gibs_78_io_ipinSE_0),
    .io_opinSE_0(gibs_78_io_opinSE_0),
    .io_ipinSW_0(gibs_78_io_ipinSW_0),
    .io_opinSW_0(gibs_78_io_opinSW_0),
    .io_itrackW_0(gibs_78_io_itrackW_0),
    .io_otrackW_0(gibs_78_io_otrackW_0),
    .io_itrackN_0(gibs_78_io_itrackN_0),
    .io_otrackN_0(gibs_78_io_otrackN_0),
    .io_itrackE_0(gibs_78_io_itrackE_0),
    .io_otrackE_0(gibs_78_io_otrackE_0)
  );
  GIB_79 gibs_79 ( // @[CGRA.scala 273:21]
    .clock(gibs_79_clock),
    .reset(gibs_79_reset),
    .io_cfg_en(gibs_79_io_cfg_en),
    .io_cfg_addr(gibs_79_io_cfg_addr),
    .io_cfg_data(gibs_79_io_cfg_data),
    .io_ipinNW_0(gibs_79_io_ipinNW_0),
    .io_ipinNW_1(gibs_79_io_ipinNW_1),
    .io_opinNW_0(gibs_79_io_opinNW_0),
    .io_ipinNE_0(gibs_79_io_ipinNE_0),
    .io_ipinNE_1(gibs_79_io_ipinNE_1),
    .io_opinNE_0(gibs_79_io_opinNE_0),
    .io_ipinSE_0(gibs_79_io_ipinSE_0),
    .io_opinSE_0(gibs_79_io_opinSE_0),
    .io_ipinSW_0(gibs_79_io_ipinSW_0),
    .io_opinSW_0(gibs_79_io_opinSW_0),
    .io_itrackW_0(gibs_79_io_itrackW_0),
    .io_otrackW_0(gibs_79_io_otrackW_0),
    .io_itrackN_0(gibs_79_io_itrackN_0),
    .io_otrackN_0(gibs_79_io_otrackN_0),
    .io_itrackE_0(gibs_79_io_itrackE_0),
    .io_otrackE_0(gibs_79_io_otrackE_0)
  );
  GIB_80 gibs_80 ( // @[CGRA.scala 273:21]
    .clock(gibs_80_clock),
    .reset(gibs_80_reset),
    .io_cfg_en(gibs_80_io_cfg_en),
    .io_cfg_addr(gibs_80_io_cfg_addr),
    .io_cfg_data(gibs_80_io_cfg_data),
    .io_ipinNW_0(gibs_80_io_ipinNW_0),
    .io_ipinNW_1(gibs_80_io_ipinNW_1),
    .io_opinNW_0(gibs_80_io_opinNW_0),
    .io_ipinSW_0(gibs_80_io_ipinSW_0),
    .io_opinSW_0(gibs_80_io_opinSW_0),
    .io_itrackW_0(gibs_80_io_itrackW_0),
    .io_otrackW_0(gibs_80_io_otrackW_0),
    .io_itrackN_0(gibs_80_io_itrackN_0),
    .io_otrackN_0(gibs_80_io_otrackN_0)
  );
  assign io_out_0 = obs_0_io_out_0; // @[CGRA.scala 345:15]
  assign io_out_1 = obs_1_io_out_0; // @[CGRA.scala 345:15]
  assign io_out_2 = obs_2_io_out_0; // @[CGRA.scala 345:15]
  assign io_out_3 = obs_3_io_out_0; // @[CGRA.scala 345:15]
  assign io_out_4 = obs_4_io_out_0; // @[CGRA.scala 345:15]
  assign io_out_5 = obs_5_io_out_0; // @[CGRA.scala 345:15]
  assign io_out_6 = obs_6_io_out_0; // @[CGRA.scala 345:15]
  assign io_out_7 = obs_7_io_out_0; // @[CGRA.scala 345:15]
  assign io_out_8 = obs_8_io_out_0; // @[CGRA.scala 345:15]
  assign io_out_9 = obs_9_io_out_0; // @[CGRA.scala 345:15]
  assign io_out_10 = obs_10_io_out_0; // @[CGRA.scala 345:15]
  assign io_out_11 = obs_11_io_out_0; // @[CGRA.scala 345:15]
  assign io_out_12 = obs_12_io_out_0; // @[CGRA.scala 345:15]
  assign io_out_13 = obs_13_io_out_0; // @[CGRA.scala 345:15]
  assign io_out_14 = obs_14_io_out_0; // @[CGRA.scala 345:15]
  assign io_out_15 = obs_15_io_out_0; // @[CGRA.scala 345:15]
  assign ibs_0_io_in_0 = io_in_0; // @[CGRA.scala 321:17]
  assign ibs_1_io_in_0 = io_in_1; // @[CGRA.scala 321:17]
  assign ibs_2_io_in_0 = io_in_2; // @[CGRA.scala 321:17]
  assign ibs_3_io_in_0 = io_in_3; // @[CGRA.scala 321:17]
  assign ibs_4_io_in_0 = io_in_4; // @[CGRA.scala 321:17]
  assign ibs_5_io_in_0 = io_in_5; // @[CGRA.scala 321:17]
  assign ibs_6_io_in_0 = io_in_6; // @[CGRA.scala 321:17]
  assign ibs_7_io_in_0 = io_in_7; // @[CGRA.scala 321:17]
  assign ibs_8_io_in_0 = io_in_8; // @[CGRA.scala 321:17]
  assign ibs_9_io_in_0 = io_in_9; // @[CGRA.scala 321:17]
  assign ibs_10_io_in_0 = io_in_10; // @[CGRA.scala 321:17]
  assign ibs_11_io_in_0 = io_in_11; // @[CGRA.scala 321:17]
  assign ibs_12_io_in_0 = io_in_12; // @[CGRA.scala 321:17]
  assign ibs_13_io_in_0 = io_in_13; // @[CGRA.scala 321:17]
  assign ibs_14_io_in_0 = io_in_14; // @[CGRA.scala 321:17]
  assign ibs_15_io_in_0 = io_in_15; // @[CGRA.scala 321:17]
  assign obs_0_clock = clock;
  assign obs_0_reset = reset;
  assign obs_0_io_cfg_en = cfgRegs_0[44]; // @[CGRA.scala 494:24]
  assign obs_0_io_cfg_addr = cfgRegs_0[43:32]; // @[CGRA.scala 495:24]
  assign obs_0_io_cfg_data = cfgRegs_0[31:0]; // @[CGRA.scala 496:24]
  assign obs_0_io_in_0 = gibs_0_io_ipinNE_0; // @[CGRA.scala 351:14]
  assign obs_0_io_in_1 = gibs_1_io_ipinNW_0; // @[CGRA.scala 355:14]
  assign obs_1_clock = clock;
  assign obs_1_reset = reset;
  assign obs_1_io_cfg_en = cfgRegs_0[44]; // @[CGRA.scala 494:24]
  assign obs_1_io_cfg_addr = cfgRegs_0[43:32]; // @[CGRA.scala 495:24]
  assign obs_1_io_cfg_data = cfgRegs_0[31:0]; // @[CGRA.scala 496:24]
  assign obs_1_io_in_0 = gibs_1_io_ipinNE_0; // @[CGRA.scala 351:14]
  assign obs_1_io_in_1 = gibs_2_io_ipinNW_0; // @[CGRA.scala 355:14]
  assign obs_2_clock = clock;
  assign obs_2_reset = reset;
  assign obs_2_io_cfg_en = cfgRegs_0[44]; // @[CGRA.scala 494:24]
  assign obs_2_io_cfg_addr = cfgRegs_0[43:32]; // @[CGRA.scala 495:24]
  assign obs_2_io_cfg_data = cfgRegs_0[31:0]; // @[CGRA.scala 496:24]
  assign obs_2_io_in_0 = gibs_2_io_ipinNE_0; // @[CGRA.scala 351:14]
  assign obs_2_io_in_1 = gibs_3_io_ipinNW_0; // @[CGRA.scala 355:14]
  assign obs_3_clock = clock;
  assign obs_3_reset = reset;
  assign obs_3_io_cfg_en = cfgRegs_0[44]; // @[CGRA.scala 494:24]
  assign obs_3_io_cfg_addr = cfgRegs_0[43:32]; // @[CGRA.scala 495:24]
  assign obs_3_io_cfg_data = cfgRegs_0[31:0]; // @[CGRA.scala 496:24]
  assign obs_3_io_in_0 = gibs_3_io_ipinNE_0; // @[CGRA.scala 351:14]
  assign obs_3_io_in_1 = gibs_4_io_ipinNW_0; // @[CGRA.scala 355:14]
  assign obs_4_clock = clock;
  assign obs_4_reset = reset;
  assign obs_4_io_cfg_en = cfgRegs_0[44]; // @[CGRA.scala 494:24]
  assign obs_4_io_cfg_addr = cfgRegs_0[43:32]; // @[CGRA.scala 495:24]
  assign obs_4_io_cfg_data = cfgRegs_0[31:0]; // @[CGRA.scala 496:24]
  assign obs_4_io_in_0 = gibs_4_io_ipinNE_0; // @[CGRA.scala 351:14]
  assign obs_4_io_in_1 = gibs_5_io_ipinNW_0; // @[CGRA.scala 355:14]
  assign obs_5_clock = clock;
  assign obs_5_reset = reset;
  assign obs_5_io_cfg_en = cfgRegs_0[44]; // @[CGRA.scala 494:24]
  assign obs_5_io_cfg_addr = cfgRegs_0[43:32]; // @[CGRA.scala 495:24]
  assign obs_5_io_cfg_data = cfgRegs_0[31:0]; // @[CGRA.scala 496:24]
  assign obs_5_io_in_0 = gibs_5_io_ipinNE_0; // @[CGRA.scala 351:14]
  assign obs_5_io_in_1 = gibs_6_io_ipinNW_0; // @[CGRA.scala 355:14]
  assign obs_6_clock = clock;
  assign obs_6_reset = reset;
  assign obs_6_io_cfg_en = cfgRegs_0[44]; // @[CGRA.scala 494:24]
  assign obs_6_io_cfg_addr = cfgRegs_0[43:32]; // @[CGRA.scala 495:24]
  assign obs_6_io_cfg_data = cfgRegs_0[31:0]; // @[CGRA.scala 496:24]
  assign obs_6_io_in_0 = gibs_6_io_ipinNE_0; // @[CGRA.scala 351:14]
  assign obs_6_io_in_1 = gibs_7_io_ipinNW_0; // @[CGRA.scala 355:14]
  assign obs_7_clock = clock;
  assign obs_7_reset = reset;
  assign obs_7_io_cfg_en = cfgRegs_0[44]; // @[CGRA.scala 494:24]
  assign obs_7_io_cfg_addr = cfgRegs_0[43:32]; // @[CGRA.scala 495:24]
  assign obs_7_io_cfg_data = cfgRegs_0[31:0]; // @[CGRA.scala 496:24]
  assign obs_7_io_in_0 = gibs_7_io_ipinNE_0; // @[CGRA.scala 351:14]
  assign obs_7_io_in_1 = gibs_8_io_ipinNW_0; // @[CGRA.scala 355:14]
  assign obs_8_clock = clock;
  assign obs_8_reset = reset;
  assign obs_8_io_cfg_en = cfgRegs_19[44]; // @[CGRA.scala 503:26]
  assign obs_8_io_cfg_addr = cfgRegs_19[43:32]; // @[CGRA.scala 504:26]
  assign obs_8_io_cfg_data = cfgRegs_19[31:0]; // @[CGRA.scala 505:26]
  assign obs_8_io_in_0 = gibs_72_io_ipinSE_0; // @[CGRA.scala 362:14]
  assign obs_8_io_in_1 = gibs_73_io_ipinSW_0; // @[CGRA.scala 366:14]
  assign obs_9_clock = clock;
  assign obs_9_reset = reset;
  assign obs_9_io_cfg_en = cfgRegs_19[44]; // @[CGRA.scala 503:26]
  assign obs_9_io_cfg_addr = cfgRegs_19[43:32]; // @[CGRA.scala 504:26]
  assign obs_9_io_cfg_data = cfgRegs_19[31:0]; // @[CGRA.scala 505:26]
  assign obs_9_io_in_0 = gibs_73_io_ipinSE_0; // @[CGRA.scala 362:14]
  assign obs_9_io_in_1 = gibs_74_io_ipinSW_0; // @[CGRA.scala 366:14]
  assign obs_10_clock = clock;
  assign obs_10_reset = reset;
  assign obs_10_io_cfg_en = cfgRegs_19[44]; // @[CGRA.scala 503:26]
  assign obs_10_io_cfg_addr = cfgRegs_19[43:32]; // @[CGRA.scala 504:26]
  assign obs_10_io_cfg_data = cfgRegs_19[31:0]; // @[CGRA.scala 505:26]
  assign obs_10_io_in_0 = gibs_74_io_ipinSE_0; // @[CGRA.scala 362:14]
  assign obs_10_io_in_1 = gibs_75_io_ipinSW_0; // @[CGRA.scala 366:14]
  assign obs_11_clock = clock;
  assign obs_11_reset = reset;
  assign obs_11_io_cfg_en = cfgRegs_19[44]; // @[CGRA.scala 503:26]
  assign obs_11_io_cfg_addr = cfgRegs_19[43:32]; // @[CGRA.scala 504:26]
  assign obs_11_io_cfg_data = cfgRegs_19[31:0]; // @[CGRA.scala 505:26]
  assign obs_11_io_in_0 = gibs_75_io_ipinSE_0; // @[CGRA.scala 362:14]
  assign obs_11_io_in_1 = gibs_76_io_ipinSW_0; // @[CGRA.scala 366:14]
  assign obs_12_clock = clock;
  assign obs_12_reset = reset;
  assign obs_12_io_cfg_en = cfgRegs_19[44]; // @[CGRA.scala 503:26]
  assign obs_12_io_cfg_addr = cfgRegs_19[43:32]; // @[CGRA.scala 504:26]
  assign obs_12_io_cfg_data = cfgRegs_19[31:0]; // @[CGRA.scala 505:26]
  assign obs_12_io_in_0 = gibs_76_io_ipinSE_0; // @[CGRA.scala 362:14]
  assign obs_12_io_in_1 = gibs_77_io_ipinSW_0; // @[CGRA.scala 366:14]
  assign obs_13_clock = clock;
  assign obs_13_reset = reset;
  assign obs_13_io_cfg_en = cfgRegs_19[44]; // @[CGRA.scala 503:26]
  assign obs_13_io_cfg_addr = cfgRegs_19[43:32]; // @[CGRA.scala 504:26]
  assign obs_13_io_cfg_data = cfgRegs_19[31:0]; // @[CGRA.scala 505:26]
  assign obs_13_io_in_0 = gibs_77_io_ipinSE_0; // @[CGRA.scala 362:14]
  assign obs_13_io_in_1 = gibs_78_io_ipinSW_0; // @[CGRA.scala 366:14]
  assign obs_14_clock = clock;
  assign obs_14_reset = reset;
  assign obs_14_io_cfg_en = cfgRegs_19[44]; // @[CGRA.scala 503:26]
  assign obs_14_io_cfg_addr = cfgRegs_19[43:32]; // @[CGRA.scala 504:26]
  assign obs_14_io_cfg_data = cfgRegs_19[31:0]; // @[CGRA.scala 505:26]
  assign obs_14_io_in_0 = gibs_78_io_ipinSE_0; // @[CGRA.scala 362:14]
  assign obs_14_io_in_1 = gibs_79_io_ipinSW_0; // @[CGRA.scala 366:14]
  assign obs_15_clock = clock;
  assign obs_15_reset = reset;
  assign obs_15_io_cfg_en = cfgRegs_19[44]; // @[CGRA.scala 503:26]
  assign obs_15_io_cfg_addr = cfgRegs_19[43:32]; // @[CGRA.scala 504:26]
  assign obs_15_io_cfg_data = cfgRegs_19[31:0]; // @[CGRA.scala 505:26]
  assign obs_15_io_in_0 = gibs_79_io_ipinSE_0; // @[CGRA.scala 362:14]
  assign obs_15_io_in_1 = gibs_80_io_ipinSW_0; // @[CGRA.scala 366:14]
  assign pes_0_clock = clock;
  assign pes_0_reset = reset;
  assign pes_0_io_cfg_en = cfgRegs_2[44]; // @[CGRA.scala 513:35]
  assign pes_0_io_cfg_addr = cfgRegs_2[43:32]; // @[CGRA.scala 514:35]
  assign pes_0_io_cfg_data = cfgRegs_2[31:0]; // @[CGRA.scala 515:35]
  assign pes_0_io_en = io_en_0; // @[CGRA.scala 377:27]
  assign pes_0_io_in_0 = gibs_0_io_ipinSE_0; // @[CGRA.scala 380:14]
  assign pes_0_io_in_1 = gibs_1_io_ipinSW_0; // @[CGRA.scala 384:14]
  assign pes_0_io_in_2 = gibs_9_io_ipinNE_0; // @[CGRA.scala 388:14]
  assign pes_0_io_in_3 = gibs_10_io_ipinNW_0; // @[CGRA.scala 392:14]
  assign pes_0_io_in_4 = gibs_0_io_ipinSE_1; // @[CGRA.scala 380:14]
  assign pes_0_io_in_5 = gibs_1_io_ipinSW_1; // @[CGRA.scala 384:14]
  assign pes_0_io_in_6 = gibs_9_io_ipinNE_1; // @[CGRA.scala 388:14]
  assign pes_0_io_in_7 = gibs_10_io_ipinNW_1; // @[CGRA.scala 392:14]
  assign pes_1_clock = clock;
  assign pes_1_reset = reset;
  assign pes_1_io_cfg_en = cfgRegs_2[44]; // @[CGRA.scala 513:35]
  assign pes_1_io_cfg_addr = cfgRegs_2[43:32]; // @[CGRA.scala 514:35]
  assign pes_1_io_cfg_data = cfgRegs_2[31:0]; // @[CGRA.scala 515:35]
  assign pes_1_io_en = io_en_1; // @[CGRA.scala 377:27]
  assign pes_1_io_in_0 = gibs_1_io_ipinSE_0; // @[CGRA.scala 380:14]
  assign pes_1_io_in_1 = gibs_2_io_ipinSW_0; // @[CGRA.scala 384:14]
  assign pes_1_io_in_2 = gibs_10_io_ipinNE_0; // @[CGRA.scala 388:14]
  assign pes_1_io_in_3 = gibs_11_io_ipinNW_0; // @[CGRA.scala 392:14]
  assign pes_1_io_in_4 = gibs_1_io_ipinSE_1; // @[CGRA.scala 380:14]
  assign pes_1_io_in_5 = gibs_2_io_ipinSW_1; // @[CGRA.scala 384:14]
  assign pes_1_io_in_6 = gibs_10_io_ipinNE_1; // @[CGRA.scala 388:14]
  assign pes_1_io_in_7 = gibs_11_io_ipinNW_1; // @[CGRA.scala 392:14]
  assign pes_2_clock = clock;
  assign pes_2_reset = reset;
  assign pes_2_io_cfg_en = cfgRegs_2[44]; // @[CGRA.scala 513:35]
  assign pes_2_io_cfg_addr = cfgRegs_2[43:32]; // @[CGRA.scala 514:35]
  assign pes_2_io_cfg_data = cfgRegs_2[31:0]; // @[CGRA.scala 515:35]
  assign pes_2_io_en = io_en_2; // @[CGRA.scala 377:27]
  assign pes_2_io_in_0 = gibs_2_io_ipinSE_0; // @[CGRA.scala 380:14]
  assign pes_2_io_in_1 = gibs_3_io_ipinSW_0; // @[CGRA.scala 384:14]
  assign pes_2_io_in_2 = gibs_11_io_ipinNE_0; // @[CGRA.scala 388:14]
  assign pes_2_io_in_3 = gibs_12_io_ipinNW_0; // @[CGRA.scala 392:14]
  assign pes_2_io_in_4 = gibs_2_io_ipinSE_1; // @[CGRA.scala 380:14]
  assign pes_2_io_in_5 = gibs_3_io_ipinSW_1; // @[CGRA.scala 384:14]
  assign pes_2_io_in_6 = gibs_11_io_ipinNE_1; // @[CGRA.scala 388:14]
  assign pes_2_io_in_7 = gibs_12_io_ipinNW_1; // @[CGRA.scala 392:14]
  assign pes_3_clock = clock;
  assign pes_3_reset = reset;
  assign pes_3_io_cfg_en = cfgRegs_2[44]; // @[CGRA.scala 513:35]
  assign pes_3_io_cfg_addr = cfgRegs_2[43:32]; // @[CGRA.scala 514:35]
  assign pes_3_io_cfg_data = cfgRegs_2[31:0]; // @[CGRA.scala 515:35]
  assign pes_3_io_en = io_en_3; // @[CGRA.scala 377:27]
  assign pes_3_io_in_0 = gibs_3_io_ipinSE_0; // @[CGRA.scala 380:14]
  assign pes_3_io_in_1 = gibs_4_io_ipinSW_0; // @[CGRA.scala 384:14]
  assign pes_3_io_in_2 = gibs_12_io_ipinNE_0; // @[CGRA.scala 388:14]
  assign pes_3_io_in_3 = gibs_13_io_ipinNW_0; // @[CGRA.scala 392:14]
  assign pes_3_io_in_4 = gibs_3_io_ipinSE_1; // @[CGRA.scala 380:14]
  assign pes_3_io_in_5 = gibs_4_io_ipinSW_1; // @[CGRA.scala 384:14]
  assign pes_3_io_in_6 = gibs_12_io_ipinNE_1; // @[CGRA.scala 388:14]
  assign pes_3_io_in_7 = gibs_13_io_ipinNW_1; // @[CGRA.scala 392:14]
  assign pes_4_clock = clock;
  assign pes_4_reset = reset;
  assign pes_4_io_cfg_en = cfgRegs_2[44]; // @[CGRA.scala 513:35]
  assign pes_4_io_cfg_addr = cfgRegs_2[43:32]; // @[CGRA.scala 514:35]
  assign pes_4_io_cfg_data = cfgRegs_2[31:0]; // @[CGRA.scala 515:35]
  assign pes_4_io_en = io_en_4; // @[CGRA.scala 377:27]
  assign pes_4_io_in_0 = gibs_4_io_ipinSE_0; // @[CGRA.scala 380:14]
  assign pes_4_io_in_1 = gibs_5_io_ipinSW_0; // @[CGRA.scala 384:14]
  assign pes_4_io_in_2 = gibs_13_io_ipinNE_0; // @[CGRA.scala 388:14]
  assign pes_4_io_in_3 = gibs_14_io_ipinNW_0; // @[CGRA.scala 392:14]
  assign pes_4_io_in_4 = gibs_4_io_ipinSE_1; // @[CGRA.scala 380:14]
  assign pes_4_io_in_5 = gibs_5_io_ipinSW_1; // @[CGRA.scala 384:14]
  assign pes_4_io_in_6 = gibs_13_io_ipinNE_1; // @[CGRA.scala 388:14]
  assign pes_4_io_in_7 = gibs_14_io_ipinNW_1; // @[CGRA.scala 392:14]
  assign pes_5_clock = clock;
  assign pes_5_reset = reset;
  assign pes_5_io_cfg_en = cfgRegs_2[44]; // @[CGRA.scala 513:35]
  assign pes_5_io_cfg_addr = cfgRegs_2[43:32]; // @[CGRA.scala 514:35]
  assign pes_5_io_cfg_data = cfgRegs_2[31:0]; // @[CGRA.scala 515:35]
  assign pes_5_io_en = io_en_5; // @[CGRA.scala 377:27]
  assign pes_5_io_in_0 = gibs_5_io_ipinSE_0; // @[CGRA.scala 380:14]
  assign pes_5_io_in_1 = gibs_6_io_ipinSW_0; // @[CGRA.scala 384:14]
  assign pes_5_io_in_2 = gibs_14_io_ipinNE_0; // @[CGRA.scala 388:14]
  assign pes_5_io_in_3 = gibs_15_io_ipinNW_0; // @[CGRA.scala 392:14]
  assign pes_5_io_in_4 = gibs_5_io_ipinSE_1; // @[CGRA.scala 380:14]
  assign pes_5_io_in_5 = gibs_6_io_ipinSW_1; // @[CGRA.scala 384:14]
  assign pes_5_io_in_6 = gibs_14_io_ipinNE_1; // @[CGRA.scala 388:14]
  assign pes_5_io_in_7 = gibs_15_io_ipinNW_1; // @[CGRA.scala 392:14]
  assign pes_6_clock = clock;
  assign pes_6_reset = reset;
  assign pes_6_io_cfg_en = cfgRegs_2[44]; // @[CGRA.scala 513:35]
  assign pes_6_io_cfg_addr = cfgRegs_2[43:32]; // @[CGRA.scala 514:35]
  assign pes_6_io_cfg_data = cfgRegs_2[31:0]; // @[CGRA.scala 515:35]
  assign pes_6_io_en = io_en_6; // @[CGRA.scala 377:27]
  assign pes_6_io_in_0 = gibs_6_io_ipinSE_0; // @[CGRA.scala 380:14]
  assign pes_6_io_in_1 = gibs_7_io_ipinSW_0; // @[CGRA.scala 384:14]
  assign pes_6_io_in_2 = gibs_15_io_ipinNE_0; // @[CGRA.scala 388:14]
  assign pes_6_io_in_3 = gibs_16_io_ipinNW_0; // @[CGRA.scala 392:14]
  assign pes_6_io_in_4 = gibs_6_io_ipinSE_1; // @[CGRA.scala 380:14]
  assign pes_6_io_in_5 = gibs_7_io_ipinSW_1; // @[CGRA.scala 384:14]
  assign pes_6_io_in_6 = gibs_15_io_ipinNE_1; // @[CGRA.scala 388:14]
  assign pes_6_io_in_7 = gibs_16_io_ipinNW_1; // @[CGRA.scala 392:14]
  assign pes_7_clock = clock;
  assign pes_7_reset = reset;
  assign pes_7_io_cfg_en = cfgRegs_2[44]; // @[CGRA.scala 513:35]
  assign pes_7_io_cfg_addr = cfgRegs_2[43:32]; // @[CGRA.scala 514:35]
  assign pes_7_io_cfg_data = cfgRegs_2[31:0]; // @[CGRA.scala 515:35]
  assign pes_7_io_en = io_en_7; // @[CGRA.scala 377:27]
  assign pes_7_io_in_0 = gibs_7_io_ipinSE_0; // @[CGRA.scala 380:14]
  assign pes_7_io_in_1 = gibs_8_io_ipinSW_0; // @[CGRA.scala 384:14]
  assign pes_7_io_in_2 = gibs_16_io_ipinNE_0; // @[CGRA.scala 388:14]
  assign pes_7_io_in_3 = gibs_17_io_ipinNW_0; // @[CGRA.scala 392:14]
  assign pes_7_io_in_4 = gibs_7_io_ipinSE_1; // @[CGRA.scala 380:14]
  assign pes_7_io_in_5 = gibs_8_io_ipinSW_1; // @[CGRA.scala 384:14]
  assign pes_7_io_in_6 = gibs_16_io_ipinNE_1; // @[CGRA.scala 388:14]
  assign pes_7_io_in_7 = gibs_17_io_ipinNW_1; // @[CGRA.scala 392:14]
  assign pes_8_clock = clock;
  assign pes_8_reset = reset;
  assign pes_8_io_cfg_en = cfgRegs_4[44]; // @[CGRA.scala 513:35]
  assign pes_8_io_cfg_addr = cfgRegs_4[43:32]; // @[CGRA.scala 514:35]
  assign pes_8_io_cfg_data = cfgRegs_4[31:0]; // @[CGRA.scala 515:35]
  assign pes_8_io_en = io_en_0; // @[CGRA.scala 377:27]
  assign pes_8_io_in_0 = gibs_9_io_ipinSE_0; // @[CGRA.scala 380:14]
  assign pes_8_io_in_1 = gibs_10_io_ipinSW_0; // @[CGRA.scala 384:14]
  assign pes_8_io_in_2 = gibs_18_io_ipinNE_0; // @[CGRA.scala 388:14]
  assign pes_8_io_in_3 = gibs_19_io_ipinNW_0; // @[CGRA.scala 392:14]
  assign pes_8_io_in_4 = gibs_9_io_ipinSE_1; // @[CGRA.scala 380:14]
  assign pes_8_io_in_5 = gibs_10_io_ipinSW_1; // @[CGRA.scala 384:14]
  assign pes_8_io_in_6 = gibs_18_io_ipinNE_1; // @[CGRA.scala 388:14]
  assign pes_8_io_in_7 = gibs_19_io_ipinNW_1; // @[CGRA.scala 392:14]
  assign pes_9_clock = clock;
  assign pes_9_reset = reset;
  assign pes_9_io_cfg_en = cfgRegs_4[44]; // @[CGRA.scala 513:35]
  assign pes_9_io_cfg_addr = cfgRegs_4[43:32]; // @[CGRA.scala 514:35]
  assign pes_9_io_cfg_data = cfgRegs_4[31:0]; // @[CGRA.scala 515:35]
  assign pes_9_io_en = io_en_1; // @[CGRA.scala 377:27]
  assign pes_9_io_in_0 = gibs_10_io_ipinSE_0; // @[CGRA.scala 380:14]
  assign pes_9_io_in_1 = gibs_11_io_ipinSW_0; // @[CGRA.scala 384:14]
  assign pes_9_io_in_2 = gibs_19_io_ipinNE_0; // @[CGRA.scala 388:14]
  assign pes_9_io_in_3 = gibs_20_io_ipinNW_0; // @[CGRA.scala 392:14]
  assign pes_9_io_in_4 = gibs_10_io_ipinSE_1; // @[CGRA.scala 380:14]
  assign pes_9_io_in_5 = gibs_11_io_ipinSW_1; // @[CGRA.scala 384:14]
  assign pes_9_io_in_6 = gibs_19_io_ipinNE_1; // @[CGRA.scala 388:14]
  assign pes_9_io_in_7 = gibs_20_io_ipinNW_1; // @[CGRA.scala 392:14]
  assign pes_10_clock = clock;
  assign pes_10_reset = reset;
  assign pes_10_io_cfg_en = cfgRegs_4[44]; // @[CGRA.scala 513:35]
  assign pes_10_io_cfg_addr = cfgRegs_4[43:32]; // @[CGRA.scala 514:35]
  assign pes_10_io_cfg_data = cfgRegs_4[31:0]; // @[CGRA.scala 515:35]
  assign pes_10_io_en = io_en_2; // @[CGRA.scala 377:27]
  assign pes_10_io_in_0 = gibs_11_io_ipinSE_0; // @[CGRA.scala 380:14]
  assign pes_10_io_in_1 = gibs_12_io_ipinSW_0; // @[CGRA.scala 384:14]
  assign pes_10_io_in_2 = gibs_20_io_ipinNE_0; // @[CGRA.scala 388:14]
  assign pes_10_io_in_3 = gibs_21_io_ipinNW_0; // @[CGRA.scala 392:14]
  assign pes_10_io_in_4 = gibs_11_io_ipinSE_1; // @[CGRA.scala 380:14]
  assign pes_10_io_in_5 = gibs_12_io_ipinSW_1; // @[CGRA.scala 384:14]
  assign pes_10_io_in_6 = gibs_20_io_ipinNE_1; // @[CGRA.scala 388:14]
  assign pes_10_io_in_7 = gibs_21_io_ipinNW_1; // @[CGRA.scala 392:14]
  assign pes_11_clock = clock;
  assign pes_11_reset = reset;
  assign pes_11_io_cfg_en = cfgRegs_4[44]; // @[CGRA.scala 513:35]
  assign pes_11_io_cfg_addr = cfgRegs_4[43:32]; // @[CGRA.scala 514:35]
  assign pes_11_io_cfg_data = cfgRegs_4[31:0]; // @[CGRA.scala 515:35]
  assign pes_11_io_en = io_en_3; // @[CGRA.scala 377:27]
  assign pes_11_io_in_0 = gibs_12_io_ipinSE_0; // @[CGRA.scala 380:14]
  assign pes_11_io_in_1 = gibs_13_io_ipinSW_0; // @[CGRA.scala 384:14]
  assign pes_11_io_in_2 = gibs_21_io_ipinNE_0; // @[CGRA.scala 388:14]
  assign pes_11_io_in_3 = gibs_22_io_ipinNW_0; // @[CGRA.scala 392:14]
  assign pes_11_io_in_4 = gibs_12_io_ipinSE_1; // @[CGRA.scala 380:14]
  assign pes_11_io_in_5 = gibs_13_io_ipinSW_1; // @[CGRA.scala 384:14]
  assign pes_11_io_in_6 = gibs_21_io_ipinNE_1; // @[CGRA.scala 388:14]
  assign pes_11_io_in_7 = gibs_22_io_ipinNW_1; // @[CGRA.scala 392:14]
  assign pes_12_clock = clock;
  assign pes_12_reset = reset;
  assign pes_12_io_cfg_en = cfgRegs_4[44]; // @[CGRA.scala 513:35]
  assign pes_12_io_cfg_addr = cfgRegs_4[43:32]; // @[CGRA.scala 514:35]
  assign pes_12_io_cfg_data = cfgRegs_4[31:0]; // @[CGRA.scala 515:35]
  assign pes_12_io_en = io_en_4; // @[CGRA.scala 377:27]
  assign pes_12_io_in_0 = gibs_13_io_ipinSE_0; // @[CGRA.scala 380:14]
  assign pes_12_io_in_1 = gibs_14_io_ipinSW_0; // @[CGRA.scala 384:14]
  assign pes_12_io_in_2 = gibs_22_io_ipinNE_0; // @[CGRA.scala 388:14]
  assign pes_12_io_in_3 = gibs_23_io_ipinNW_0; // @[CGRA.scala 392:14]
  assign pes_12_io_in_4 = gibs_13_io_ipinSE_1; // @[CGRA.scala 380:14]
  assign pes_12_io_in_5 = gibs_14_io_ipinSW_1; // @[CGRA.scala 384:14]
  assign pes_12_io_in_6 = gibs_22_io_ipinNE_1; // @[CGRA.scala 388:14]
  assign pes_12_io_in_7 = gibs_23_io_ipinNW_1; // @[CGRA.scala 392:14]
  assign pes_13_clock = clock;
  assign pes_13_reset = reset;
  assign pes_13_io_cfg_en = cfgRegs_4[44]; // @[CGRA.scala 513:35]
  assign pes_13_io_cfg_addr = cfgRegs_4[43:32]; // @[CGRA.scala 514:35]
  assign pes_13_io_cfg_data = cfgRegs_4[31:0]; // @[CGRA.scala 515:35]
  assign pes_13_io_en = io_en_5; // @[CGRA.scala 377:27]
  assign pes_13_io_in_0 = gibs_14_io_ipinSE_0; // @[CGRA.scala 380:14]
  assign pes_13_io_in_1 = gibs_15_io_ipinSW_0; // @[CGRA.scala 384:14]
  assign pes_13_io_in_2 = gibs_23_io_ipinNE_0; // @[CGRA.scala 388:14]
  assign pes_13_io_in_3 = gibs_24_io_ipinNW_0; // @[CGRA.scala 392:14]
  assign pes_13_io_in_4 = gibs_14_io_ipinSE_1; // @[CGRA.scala 380:14]
  assign pes_13_io_in_5 = gibs_15_io_ipinSW_1; // @[CGRA.scala 384:14]
  assign pes_13_io_in_6 = gibs_23_io_ipinNE_1; // @[CGRA.scala 388:14]
  assign pes_13_io_in_7 = gibs_24_io_ipinNW_1; // @[CGRA.scala 392:14]
  assign pes_14_clock = clock;
  assign pes_14_reset = reset;
  assign pes_14_io_cfg_en = cfgRegs_4[44]; // @[CGRA.scala 513:35]
  assign pes_14_io_cfg_addr = cfgRegs_4[43:32]; // @[CGRA.scala 514:35]
  assign pes_14_io_cfg_data = cfgRegs_4[31:0]; // @[CGRA.scala 515:35]
  assign pes_14_io_en = io_en_6; // @[CGRA.scala 377:27]
  assign pes_14_io_in_0 = gibs_15_io_ipinSE_0; // @[CGRA.scala 380:14]
  assign pes_14_io_in_1 = gibs_16_io_ipinSW_0; // @[CGRA.scala 384:14]
  assign pes_14_io_in_2 = gibs_24_io_ipinNE_0; // @[CGRA.scala 388:14]
  assign pes_14_io_in_3 = gibs_25_io_ipinNW_0; // @[CGRA.scala 392:14]
  assign pes_14_io_in_4 = gibs_15_io_ipinSE_1; // @[CGRA.scala 380:14]
  assign pes_14_io_in_5 = gibs_16_io_ipinSW_1; // @[CGRA.scala 384:14]
  assign pes_14_io_in_6 = gibs_24_io_ipinNE_1; // @[CGRA.scala 388:14]
  assign pes_14_io_in_7 = gibs_25_io_ipinNW_1; // @[CGRA.scala 392:14]
  assign pes_15_clock = clock;
  assign pes_15_reset = reset;
  assign pes_15_io_cfg_en = cfgRegs_4[44]; // @[CGRA.scala 513:35]
  assign pes_15_io_cfg_addr = cfgRegs_4[43:32]; // @[CGRA.scala 514:35]
  assign pes_15_io_cfg_data = cfgRegs_4[31:0]; // @[CGRA.scala 515:35]
  assign pes_15_io_en = io_en_7; // @[CGRA.scala 377:27]
  assign pes_15_io_in_0 = gibs_16_io_ipinSE_0; // @[CGRA.scala 380:14]
  assign pes_15_io_in_1 = gibs_17_io_ipinSW_0; // @[CGRA.scala 384:14]
  assign pes_15_io_in_2 = gibs_25_io_ipinNE_0; // @[CGRA.scala 388:14]
  assign pes_15_io_in_3 = gibs_26_io_ipinNW_0; // @[CGRA.scala 392:14]
  assign pes_15_io_in_4 = gibs_16_io_ipinSE_1; // @[CGRA.scala 380:14]
  assign pes_15_io_in_5 = gibs_17_io_ipinSW_1; // @[CGRA.scala 384:14]
  assign pes_15_io_in_6 = gibs_25_io_ipinNE_1; // @[CGRA.scala 388:14]
  assign pes_15_io_in_7 = gibs_26_io_ipinNW_1; // @[CGRA.scala 392:14]
  assign pes_16_clock = clock;
  assign pes_16_reset = reset;
  assign pes_16_io_cfg_en = cfgRegs_6[44]; // @[CGRA.scala 513:35]
  assign pes_16_io_cfg_addr = cfgRegs_6[43:32]; // @[CGRA.scala 514:35]
  assign pes_16_io_cfg_data = cfgRegs_6[31:0]; // @[CGRA.scala 515:35]
  assign pes_16_io_en = io_en_0; // @[CGRA.scala 377:27]
  assign pes_16_io_in_0 = gibs_18_io_ipinSE_0; // @[CGRA.scala 380:14]
  assign pes_16_io_in_1 = gibs_19_io_ipinSW_0; // @[CGRA.scala 384:14]
  assign pes_16_io_in_2 = gibs_27_io_ipinNE_0; // @[CGRA.scala 388:14]
  assign pes_16_io_in_3 = gibs_28_io_ipinNW_0; // @[CGRA.scala 392:14]
  assign pes_16_io_in_4 = gibs_18_io_ipinSE_1; // @[CGRA.scala 380:14]
  assign pes_16_io_in_5 = gibs_19_io_ipinSW_1; // @[CGRA.scala 384:14]
  assign pes_16_io_in_6 = gibs_27_io_ipinNE_1; // @[CGRA.scala 388:14]
  assign pes_16_io_in_7 = gibs_28_io_ipinNW_1; // @[CGRA.scala 392:14]
  assign pes_17_clock = clock;
  assign pes_17_reset = reset;
  assign pes_17_io_cfg_en = cfgRegs_6[44]; // @[CGRA.scala 513:35]
  assign pes_17_io_cfg_addr = cfgRegs_6[43:32]; // @[CGRA.scala 514:35]
  assign pes_17_io_cfg_data = cfgRegs_6[31:0]; // @[CGRA.scala 515:35]
  assign pes_17_io_en = io_en_1; // @[CGRA.scala 377:27]
  assign pes_17_io_in_0 = gibs_19_io_ipinSE_0; // @[CGRA.scala 380:14]
  assign pes_17_io_in_1 = gibs_20_io_ipinSW_0; // @[CGRA.scala 384:14]
  assign pes_17_io_in_2 = gibs_28_io_ipinNE_0; // @[CGRA.scala 388:14]
  assign pes_17_io_in_3 = gibs_29_io_ipinNW_0; // @[CGRA.scala 392:14]
  assign pes_17_io_in_4 = gibs_19_io_ipinSE_1; // @[CGRA.scala 380:14]
  assign pes_17_io_in_5 = gibs_20_io_ipinSW_1; // @[CGRA.scala 384:14]
  assign pes_17_io_in_6 = gibs_28_io_ipinNE_1; // @[CGRA.scala 388:14]
  assign pes_17_io_in_7 = gibs_29_io_ipinNW_1; // @[CGRA.scala 392:14]
  assign pes_18_clock = clock;
  assign pes_18_reset = reset;
  assign pes_18_io_cfg_en = cfgRegs_6[44]; // @[CGRA.scala 513:35]
  assign pes_18_io_cfg_addr = cfgRegs_6[43:32]; // @[CGRA.scala 514:35]
  assign pes_18_io_cfg_data = cfgRegs_6[31:0]; // @[CGRA.scala 515:35]
  assign pes_18_io_en = io_en_2; // @[CGRA.scala 377:27]
  assign pes_18_io_in_0 = gibs_20_io_ipinSE_0; // @[CGRA.scala 380:14]
  assign pes_18_io_in_1 = gibs_21_io_ipinSW_0; // @[CGRA.scala 384:14]
  assign pes_18_io_in_2 = gibs_29_io_ipinNE_0; // @[CGRA.scala 388:14]
  assign pes_18_io_in_3 = gibs_30_io_ipinNW_0; // @[CGRA.scala 392:14]
  assign pes_18_io_in_4 = gibs_20_io_ipinSE_1; // @[CGRA.scala 380:14]
  assign pes_18_io_in_5 = gibs_21_io_ipinSW_1; // @[CGRA.scala 384:14]
  assign pes_18_io_in_6 = gibs_29_io_ipinNE_1; // @[CGRA.scala 388:14]
  assign pes_18_io_in_7 = gibs_30_io_ipinNW_1; // @[CGRA.scala 392:14]
  assign pes_19_clock = clock;
  assign pes_19_reset = reset;
  assign pes_19_io_cfg_en = cfgRegs_6[44]; // @[CGRA.scala 513:35]
  assign pes_19_io_cfg_addr = cfgRegs_6[43:32]; // @[CGRA.scala 514:35]
  assign pes_19_io_cfg_data = cfgRegs_6[31:0]; // @[CGRA.scala 515:35]
  assign pes_19_io_en = io_en_3; // @[CGRA.scala 377:27]
  assign pes_19_io_in_0 = gibs_21_io_ipinSE_0; // @[CGRA.scala 380:14]
  assign pes_19_io_in_1 = gibs_22_io_ipinSW_0; // @[CGRA.scala 384:14]
  assign pes_19_io_in_2 = gibs_30_io_ipinNE_0; // @[CGRA.scala 388:14]
  assign pes_19_io_in_3 = gibs_31_io_ipinNW_0; // @[CGRA.scala 392:14]
  assign pes_19_io_in_4 = gibs_21_io_ipinSE_1; // @[CGRA.scala 380:14]
  assign pes_19_io_in_5 = gibs_22_io_ipinSW_1; // @[CGRA.scala 384:14]
  assign pes_19_io_in_6 = gibs_30_io_ipinNE_1; // @[CGRA.scala 388:14]
  assign pes_19_io_in_7 = gibs_31_io_ipinNW_1; // @[CGRA.scala 392:14]
  assign pes_20_clock = clock;
  assign pes_20_reset = reset;
  assign pes_20_io_cfg_en = cfgRegs_6[44]; // @[CGRA.scala 513:35]
  assign pes_20_io_cfg_addr = cfgRegs_6[43:32]; // @[CGRA.scala 514:35]
  assign pes_20_io_cfg_data = cfgRegs_6[31:0]; // @[CGRA.scala 515:35]
  assign pes_20_io_en = io_en_4; // @[CGRA.scala 377:27]
  assign pes_20_io_in_0 = gibs_22_io_ipinSE_0; // @[CGRA.scala 380:14]
  assign pes_20_io_in_1 = gibs_23_io_ipinSW_0; // @[CGRA.scala 384:14]
  assign pes_20_io_in_2 = gibs_31_io_ipinNE_0; // @[CGRA.scala 388:14]
  assign pes_20_io_in_3 = gibs_32_io_ipinNW_0; // @[CGRA.scala 392:14]
  assign pes_20_io_in_4 = gibs_22_io_ipinSE_1; // @[CGRA.scala 380:14]
  assign pes_20_io_in_5 = gibs_23_io_ipinSW_1; // @[CGRA.scala 384:14]
  assign pes_20_io_in_6 = gibs_31_io_ipinNE_1; // @[CGRA.scala 388:14]
  assign pes_20_io_in_7 = gibs_32_io_ipinNW_1; // @[CGRA.scala 392:14]
  assign pes_21_clock = clock;
  assign pes_21_reset = reset;
  assign pes_21_io_cfg_en = cfgRegs_6[44]; // @[CGRA.scala 513:35]
  assign pes_21_io_cfg_addr = cfgRegs_6[43:32]; // @[CGRA.scala 514:35]
  assign pes_21_io_cfg_data = cfgRegs_6[31:0]; // @[CGRA.scala 515:35]
  assign pes_21_io_en = io_en_5; // @[CGRA.scala 377:27]
  assign pes_21_io_in_0 = gibs_23_io_ipinSE_0; // @[CGRA.scala 380:14]
  assign pes_21_io_in_1 = gibs_24_io_ipinSW_0; // @[CGRA.scala 384:14]
  assign pes_21_io_in_2 = gibs_32_io_ipinNE_0; // @[CGRA.scala 388:14]
  assign pes_21_io_in_3 = gibs_33_io_ipinNW_0; // @[CGRA.scala 392:14]
  assign pes_21_io_in_4 = gibs_23_io_ipinSE_1; // @[CGRA.scala 380:14]
  assign pes_21_io_in_5 = gibs_24_io_ipinSW_1; // @[CGRA.scala 384:14]
  assign pes_21_io_in_6 = gibs_32_io_ipinNE_1; // @[CGRA.scala 388:14]
  assign pes_21_io_in_7 = gibs_33_io_ipinNW_1; // @[CGRA.scala 392:14]
  assign pes_22_clock = clock;
  assign pes_22_reset = reset;
  assign pes_22_io_cfg_en = cfgRegs_6[44]; // @[CGRA.scala 513:35]
  assign pes_22_io_cfg_addr = cfgRegs_6[43:32]; // @[CGRA.scala 514:35]
  assign pes_22_io_cfg_data = cfgRegs_6[31:0]; // @[CGRA.scala 515:35]
  assign pes_22_io_en = io_en_6; // @[CGRA.scala 377:27]
  assign pes_22_io_in_0 = gibs_24_io_ipinSE_0; // @[CGRA.scala 380:14]
  assign pes_22_io_in_1 = gibs_25_io_ipinSW_0; // @[CGRA.scala 384:14]
  assign pes_22_io_in_2 = gibs_33_io_ipinNE_0; // @[CGRA.scala 388:14]
  assign pes_22_io_in_3 = gibs_34_io_ipinNW_0; // @[CGRA.scala 392:14]
  assign pes_22_io_in_4 = gibs_24_io_ipinSE_1; // @[CGRA.scala 380:14]
  assign pes_22_io_in_5 = gibs_25_io_ipinSW_1; // @[CGRA.scala 384:14]
  assign pes_22_io_in_6 = gibs_33_io_ipinNE_1; // @[CGRA.scala 388:14]
  assign pes_22_io_in_7 = gibs_34_io_ipinNW_1; // @[CGRA.scala 392:14]
  assign pes_23_clock = clock;
  assign pes_23_reset = reset;
  assign pes_23_io_cfg_en = cfgRegs_6[44]; // @[CGRA.scala 513:35]
  assign pes_23_io_cfg_addr = cfgRegs_6[43:32]; // @[CGRA.scala 514:35]
  assign pes_23_io_cfg_data = cfgRegs_6[31:0]; // @[CGRA.scala 515:35]
  assign pes_23_io_en = io_en_7; // @[CGRA.scala 377:27]
  assign pes_23_io_in_0 = gibs_25_io_ipinSE_0; // @[CGRA.scala 380:14]
  assign pes_23_io_in_1 = gibs_26_io_ipinSW_0; // @[CGRA.scala 384:14]
  assign pes_23_io_in_2 = gibs_34_io_ipinNE_0; // @[CGRA.scala 388:14]
  assign pes_23_io_in_3 = gibs_35_io_ipinNW_0; // @[CGRA.scala 392:14]
  assign pes_23_io_in_4 = gibs_25_io_ipinSE_1; // @[CGRA.scala 380:14]
  assign pes_23_io_in_5 = gibs_26_io_ipinSW_1; // @[CGRA.scala 384:14]
  assign pes_23_io_in_6 = gibs_34_io_ipinNE_1; // @[CGRA.scala 388:14]
  assign pes_23_io_in_7 = gibs_35_io_ipinNW_1; // @[CGRA.scala 392:14]
  assign pes_24_clock = clock;
  assign pes_24_reset = reset;
  assign pes_24_io_cfg_en = cfgRegs_8[44]; // @[CGRA.scala 513:35]
  assign pes_24_io_cfg_addr = cfgRegs_8[43:32]; // @[CGRA.scala 514:35]
  assign pes_24_io_cfg_data = cfgRegs_8[31:0]; // @[CGRA.scala 515:35]
  assign pes_24_io_en = io_en_0; // @[CGRA.scala 377:27]
  assign pes_24_io_in_0 = gibs_27_io_ipinSE_0; // @[CGRA.scala 380:14]
  assign pes_24_io_in_1 = gibs_28_io_ipinSW_0; // @[CGRA.scala 384:14]
  assign pes_24_io_in_2 = gibs_36_io_ipinNE_0; // @[CGRA.scala 388:14]
  assign pes_24_io_in_3 = gibs_37_io_ipinNW_0; // @[CGRA.scala 392:14]
  assign pes_24_io_in_4 = gibs_27_io_ipinSE_1; // @[CGRA.scala 380:14]
  assign pes_24_io_in_5 = gibs_28_io_ipinSW_1; // @[CGRA.scala 384:14]
  assign pes_24_io_in_6 = gibs_36_io_ipinNE_1; // @[CGRA.scala 388:14]
  assign pes_24_io_in_7 = gibs_37_io_ipinNW_1; // @[CGRA.scala 392:14]
  assign pes_25_clock = clock;
  assign pes_25_reset = reset;
  assign pes_25_io_cfg_en = cfgRegs_8[44]; // @[CGRA.scala 513:35]
  assign pes_25_io_cfg_addr = cfgRegs_8[43:32]; // @[CGRA.scala 514:35]
  assign pes_25_io_cfg_data = cfgRegs_8[31:0]; // @[CGRA.scala 515:35]
  assign pes_25_io_en = io_en_1; // @[CGRA.scala 377:27]
  assign pes_25_io_in_0 = gibs_28_io_ipinSE_0; // @[CGRA.scala 380:14]
  assign pes_25_io_in_1 = gibs_29_io_ipinSW_0; // @[CGRA.scala 384:14]
  assign pes_25_io_in_2 = gibs_37_io_ipinNE_0; // @[CGRA.scala 388:14]
  assign pes_25_io_in_3 = gibs_38_io_ipinNW_0; // @[CGRA.scala 392:14]
  assign pes_25_io_in_4 = gibs_28_io_ipinSE_1; // @[CGRA.scala 380:14]
  assign pes_25_io_in_5 = gibs_29_io_ipinSW_1; // @[CGRA.scala 384:14]
  assign pes_25_io_in_6 = gibs_37_io_ipinNE_1; // @[CGRA.scala 388:14]
  assign pes_25_io_in_7 = gibs_38_io_ipinNW_1; // @[CGRA.scala 392:14]
  assign pes_26_clock = clock;
  assign pes_26_reset = reset;
  assign pes_26_io_cfg_en = cfgRegs_8[44]; // @[CGRA.scala 513:35]
  assign pes_26_io_cfg_addr = cfgRegs_8[43:32]; // @[CGRA.scala 514:35]
  assign pes_26_io_cfg_data = cfgRegs_8[31:0]; // @[CGRA.scala 515:35]
  assign pes_26_io_en = io_en_2; // @[CGRA.scala 377:27]
  assign pes_26_io_in_0 = gibs_29_io_ipinSE_0; // @[CGRA.scala 380:14]
  assign pes_26_io_in_1 = gibs_30_io_ipinSW_0; // @[CGRA.scala 384:14]
  assign pes_26_io_in_2 = gibs_38_io_ipinNE_0; // @[CGRA.scala 388:14]
  assign pes_26_io_in_3 = gibs_39_io_ipinNW_0; // @[CGRA.scala 392:14]
  assign pes_26_io_in_4 = gibs_29_io_ipinSE_1; // @[CGRA.scala 380:14]
  assign pes_26_io_in_5 = gibs_30_io_ipinSW_1; // @[CGRA.scala 384:14]
  assign pes_26_io_in_6 = gibs_38_io_ipinNE_1; // @[CGRA.scala 388:14]
  assign pes_26_io_in_7 = gibs_39_io_ipinNW_1; // @[CGRA.scala 392:14]
  assign pes_27_clock = clock;
  assign pes_27_reset = reset;
  assign pes_27_io_cfg_en = cfgRegs_8[44]; // @[CGRA.scala 513:35]
  assign pes_27_io_cfg_addr = cfgRegs_8[43:32]; // @[CGRA.scala 514:35]
  assign pes_27_io_cfg_data = cfgRegs_8[31:0]; // @[CGRA.scala 515:35]
  assign pes_27_io_en = io_en_3; // @[CGRA.scala 377:27]
  assign pes_27_io_in_0 = gibs_30_io_ipinSE_0; // @[CGRA.scala 380:14]
  assign pes_27_io_in_1 = gibs_31_io_ipinSW_0; // @[CGRA.scala 384:14]
  assign pes_27_io_in_2 = gibs_39_io_ipinNE_0; // @[CGRA.scala 388:14]
  assign pes_27_io_in_3 = gibs_40_io_ipinNW_0; // @[CGRA.scala 392:14]
  assign pes_27_io_in_4 = gibs_30_io_ipinSE_1; // @[CGRA.scala 380:14]
  assign pes_27_io_in_5 = gibs_31_io_ipinSW_1; // @[CGRA.scala 384:14]
  assign pes_27_io_in_6 = gibs_39_io_ipinNE_1; // @[CGRA.scala 388:14]
  assign pes_27_io_in_7 = gibs_40_io_ipinNW_1; // @[CGRA.scala 392:14]
  assign pes_28_clock = clock;
  assign pes_28_reset = reset;
  assign pes_28_io_cfg_en = cfgRegs_8[44]; // @[CGRA.scala 513:35]
  assign pes_28_io_cfg_addr = cfgRegs_8[43:32]; // @[CGRA.scala 514:35]
  assign pes_28_io_cfg_data = cfgRegs_8[31:0]; // @[CGRA.scala 515:35]
  assign pes_28_io_en = io_en_4; // @[CGRA.scala 377:27]
  assign pes_28_io_in_0 = gibs_31_io_ipinSE_0; // @[CGRA.scala 380:14]
  assign pes_28_io_in_1 = gibs_32_io_ipinSW_0; // @[CGRA.scala 384:14]
  assign pes_28_io_in_2 = gibs_40_io_ipinNE_0; // @[CGRA.scala 388:14]
  assign pes_28_io_in_3 = gibs_41_io_ipinNW_0; // @[CGRA.scala 392:14]
  assign pes_28_io_in_4 = gibs_31_io_ipinSE_1; // @[CGRA.scala 380:14]
  assign pes_28_io_in_5 = gibs_32_io_ipinSW_1; // @[CGRA.scala 384:14]
  assign pes_28_io_in_6 = gibs_40_io_ipinNE_1; // @[CGRA.scala 388:14]
  assign pes_28_io_in_7 = gibs_41_io_ipinNW_1; // @[CGRA.scala 392:14]
  assign pes_29_clock = clock;
  assign pes_29_reset = reset;
  assign pes_29_io_cfg_en = cfgRegs_8[44]; // @[CGRA.scala 513:35]
  assign pes_29_io_cfg_addr = cfgRegs_8[43:32]; // @[CGRA.scala 514:35]
  assign pes_29_io_cfg_data = cfgRegs_8[31:0]; // @[CGRA.scala 515:35]
  assign pes_29_io_en = io_en_5; // @[CGRA.scala 377:27]
  assign pes_29_io_in_0 = gibs_32_io_ipinSE_0; // @[CGRA.scala 380:14]
  assign pes_29_io_in_1 = gibs_33_io_ipinSW_0; // @[CGRA.scala 384:14]
  assign pes_29_io_in_2 = gibs_41_io_ipinNE_0; // @[CGRA.scala 388:14]
  assign pes_29_io_in_3 = gibs_42_io_ipinNW_0; // @[CGRA.scala 392:14]
  assign pes_29_io_in_4 = gibs_32_io_ipinSE_1; // @[CGRA.scala 380:14]
  assign pes_29_io_in_5 = gibs_33_io_ipinSW_1; // @[CGRA.scala 384:14]
  assign pes_29_io_in_6 = gibs_41_io_ipinNE_1; // @[CGRA.scala 388:14]
  assign pes_29_io_in_7 = gibs_42_io_ipinNW_1; // @[CGRA.scala 392:14]
  assign pes_30_clock = clock;
  assign pes_30_reset = reset;
  assign pes_30_io_cfg_en = cfgRegs_8[44]; // @[CGRA.scala 513:35]
  assign pes_30_io_cfg_addr = cfgRegs_8[43:32]; // @[CGRA.scala 514:35]
  assign pes_30_io_cfg_data = cfgRegs_8[31:0]; // @[CGRA.scala 515:35]
  assign pes_30_io_en = io_en_6; // @[CGRA.scala 377:27]
  assign pes_30_io_in_0 = gibs_33_io_ipinSE_0; // @[CGRA.scala 380:14]
  assign pes_30_io_in_1 = gibs_34_io_ipinSW_0; // @[CGRA.scala 384:14]
  assign pes_30_io_in_2 = gibs_42_io_ipinNE_0; // @[CGRA.scala 388:14]
  assign pes_30_io_in_3 = gibs_43_io_ipinNW_0; // @[CGRA.scala 392:14]
  assign pes_30_io_in_4 = gibs_33_io_ipinSE_1; // @[CGRA.scala 380:14]
  assign pes_30_io_in_5 = gibs_34_io_ipinSW_1; // @[CGRA.scala 384:14]
  assign pes_30_io_in_6 = gibs_42_io_ipinNE_1; // @[CGRA.scala 388:14]
  assign pes_30_io_in_7 = gibs_43_io_ipinNW_1; // @[CGRA.scala 392:14]
  assign pes_31_clock = clock;
  assign pes_31_reset = reset;
  assign pes_31_io_cfg_en = cfgRegs_8[44]; // @[CGRA.scala 513:35]
  assign pes_31_io_cfg_addr = cfgRegs_8[43:32]; // @[CGRA.scala 514:35]
  assign pes_31_io_cfg_data = cfgRegs_8[31:0]; // @[CGRA.scala 515:35]
  assign pes_31_io_en = io_en_7; // @[CGRA.scala 377:27]
  assign pes_31_io_in_0 = gibs_34_io_ipinSE_0; // @[CGRA.scala 380:14]
  assign pes_31_io_in_1 = gibs_35_io_ipinSW_0; // @[CGRA.scala 384:14]
  assign pes_31_io_in_2 = gibs_43_io_ipinNE_0; // @[CGRA.scala 388:14]
  assign pes_31_io_in_3 = gibs_44_io_ipinNW_0; // @[CGRA.scala 392:14]
  assign pes_31_io_in_4 = gibs_34_io_ipinSE_1; // @[CGRA.scala 380:14]
  assign pes_31_io_in_5 = gibs_35_io_ipinSW_1; // @[CGRA.scala 384:14]
  assign pes_31_io_in_6 = gibs_43_io_ipinNE_1; // @[CGRA.scala 388:14]
  assign pes_31_io_in_7 = gibs_44_io_ipinNW_1; // @[CGRA.scala 392:14]
  assign pes_32_clock = clock;
  assign pes_32_reset = reset;
  assign pes_32_io_cfg_en = cfgRegs_10[44]; // @[CGRA.scala 513:35]
  assign pes_32_io_cfg_addr = cfgRegs_10[43:32]; // @[CGRA.scala 514:35]
  assign pes_32_io_cfg_data = cfgRegs_10[31:0]; // @[CGRA.scala 515:35]
  assign pes_32_io_en = io_en_0; // @[CGRA.scala 377:27]
  assign pes_32_io_in_0 = gibs_36_io_ipinSE_0; // @[CGRA.scala 380:14]
  assign pes_32_io_in_1 = gibs_37_io_ipinSW_0; // @[CGRA.scala 384:14]
  assign pes_32_io_in_2 = gibs_45_io_ipinNE_0; // @[CGRA.scala 388:14]
  assign pes_32_io_in_3 = gibs_46_io_ipinNW_0; // @[CGRA.scala 392:14]
  assign pes_32_io_in_4 = gibs_36_io_ipinSE_1; // @[CGRA.scala 380:14]
  assign pes_32_io_in_5 = gibs_37_io_ipinSW_1; // @[CGRA.scala 384:14]
  assign pes_32_io_in_6 = gibs_45_io_ipinNE_1; // @[CGRA.scala 388:14]
  assign pes_32_io_in_7 = gibs_46_io_ipinNW_1; // @[CGRA.scala 392:14]
  assign pes_33_clock = clock;
  assign pes_33_reset = reset;
  assign pes_33_io_cfg_en = cfgRegs_10[44]; // @[CGRA.scala 513:35]
  assign pes_33_io_cfg_addr = cfgRegs_10[43:32]; // @[CGRA.scala 514:35]
  assign pes_33_io_cfg_data = cfgRegs_10[31:0]; // @[CGRA.scala 515:35]
  assign pes_33_io_en = io_en_1; // @[CGRA.scala 377:27]
  assign pes_33_io_in_0 = gibs_37_io_ipinSE_0; // @[CGRA.scala 380:14]
  assign pes_33_io_in_1 = gibs_38_io_ipinSW_0; // @[CGRA.scala 384:14]
  assign pes_33_io_in_2 = gibs_46_io_ipinNE_0; // @[CGRA.scala 388:14]
  assign pes_33_io_in_3 = gibs_47_io_ipinNW_0; // @[CGRA.scala 392:14]
  assign pes_33_io_in_4 = gibs_37_io_ipinSE_1; // @[CGRA.scala 380:14]
  assign pes_33_io_in_5 = gibs_38_io_ipinSW_1; // @[CGRA.scala 384:14]
  assign pes_33_io_in_6 = gibs_46_io_ipinNE_1; // @[CGRA.scala 388:14]
  assign pes_33_io_in_7 = gibs_47_io_ipinNW_1; // @[CGRA.scala 392:14]
  assign pes_34_clock = clock;
  assign pes_34_reset = reset;
  assign pes_34_io_cfg_en = cfgRegs_10[44]; // @[CGRA.scala 513:35]
  assign pes_34_io_cfg_addr = cfgRegs_10[43:32]; // @[CGRA.scala 514:35]
  assign pes_34_io_cfg_data = cfgRegs_10[31:0]; // @[CGRA.scala 515:35]
  assign pes_34_io_en = io_en_2; // @[CGRA.scala 377:27]
  assign pes_34_io_in_0 = gibs_38_io_ipinSE_0; // @[CGRA.scala 380:14]
  assign pes_34_io_in_1 = gibs_39_io_ipinSW_0; // @[CGRA.scala 384:14]
  assign pes_34_io_in_2 = gibs_47_io_ipinNE_0; // @[CGRA.scala 388:14]
  assign pes_34_io_in_3 = gibs_48_io_ipinNW_0; // @[CGRA.scala 392:14]
  assign pes_34_io_in_4 = gibs_38_io_ipinSE_1; // @[CGRA.scala 380:14]
  assign pes_34_io_in_5 = gibs_39_io_ipinSW_1; // @[CGRA.scala 384:14]
  assign pes_34_io_in_6 = gibs_47_io_ipinNE_1; // @[CGRA.scala 388:14]
  assign pes_34_io_in_7 = gibs_48_io_ipinNW_1; // @[CGRA.scala 392:14]
  assign pes_35_clock = clock;
  assign pes_35_reset = reset;
  assign pes_35_io_cfg_en = cfgRegs_10[44]; // @[CGRA.scala 513:35]
  assign pes_35_io_cfg_addr = cfgRegs_10[43:32]; // @[CGRA.scala 514:35]
  assign pes_35_io_cfg_data = cfgRegs_10[31:0]; // @[CGRA.scala 515:35]
  assign pes_35_io_en = io_en_3; // @[CGRA.scala 377:27]
  assign pes_35_io_in_0 = gibs_39_io_ipinSE_0; // @[CGRA.scala 380:14]
  assign pes_35_io_in_1 = gibs_40_io_ipinSW_0; // @[CGRA.scala 384:14]
  assign pes_35_io_in_2 = gibs_48_io_ipinNE_0; // @[CGRA.scala 388:14]
  assign pes_35_io_in_3 = gibs_49_io_ipinNW_0; // @[CGRA.scala 392:14]
  assign pes_35_io_in_4 = gibs_39_io_ipinSE_1; // @[CGRA.scala 380:14]
  assign pes_35_io_in_5 = gibs_40_io_ipinSW_1; // @[CGRA.scala 384:14]
  assign pes_35_io_in_6 = gibs_48_io_ipinNE_1; // @[CGRA.scala 388:14]
  assign pes_35_io_in_7 = gibs_49_io_ipinNW_1; // @[CGRA.scala 392:14]
  assign pes_36_clock = clock;
  assign pes_36_reset = reset;
  assign pes_36_io_cfg_en = cfgRegs_10[44]; // @[CGRA.scala 513:35]
  assign pes_36_io_cfg_addr = cfgRegs_10[43:32]; // @[CGRA.scala 514:35]
  assign pes_36_io_cfg_data = cfgRegs_10[31:0]; // @[CGRA.scala 515:35]
  assign pes_36_io_en = io_en_4; // @[CGRA.scala 377:27]
  assign pes_36_io_in_0 = gibs_40_io_ipinSE_0; // @[CGRA.scala 380:14]
  assign pes_36_io_in_1 = gibs_41_io_ipinSW_0; // @[CGRA.scala 384:14]
  assign pes_36_io_in_2 = gibs_49_io_ipinNE_0; // @[CGRA.scala 388:14]
  assign pes_36_io_in_3 = gibs_50_io_ipinNW_0; // @[CGRA.scala 392:14]
  assign pes_36_io_in_4 = gibs_40_io_ipinSE_1; // @[CGRA.scala 380:14]
  assign pes_36_io_in_5 = gibs_41_io_ipinSW_1; // @[CGRA.scala 384:14]
  assign pes_36_io_in_6 = gibs_49_io_ipinNE_1; // @[CGRA.scala 388:14]
  assign pes_36_io_in_7 = gibs_50_io_ipinNW_1; // @[CGRA.scala 392:14]
  assign pes_37_clock = clock;
  assign pes_37_reset = reset;
  assign pes_37_io_cfg_en = cfgRegs_10[44]; // @[CGRA.scala 513:35]
  assign pes_37_io_cfg_addr = cfgRegs_10[43:32]; // @[CGRA.scala 514:35]
  assign pes_37_io_cfg_data = cfgRegs_10[31:0]; // @[CGRA.scala 515:35]
  assign pes_37_io_en = io_en_5; // @[CGRA.scala 377:27]
  assign pes_37_io_in_0 = gibs_41_io_ipinSE_0; // @[CGRA.scala 380:14]
  assign pes_37_io_in_1 = gibs_42_io_ipinSW_0; // @[CGRA.scala 384:14]
  assign pes_37_io_in_2 = gibs_50_io_ipinNE_0; // @[CGRA.scala 388:14]
  assign pes_37_io_in_3 = gibs_51_io_ipinNW_0; // @[CGRA.scala 392:14]
  assign pes_37_io_in_4 = gibs_41_io_ipinSE_1; // @[CGRA.scala 380:14]
  assign pes_37_io_in_5 = gibs_42_io_ipinSW_1; // @[CGRA.scala 384:14]
  assign pes_37_io_in_6 = gibs_50_io_ipinNE_1; // @[CGRA.scala 388:14]
  assign pes_37_io_in_7 = gibs_51_io_ipinNW_1; // @[CGRA.scala 392:14]
  assign pes_38_clock = clock;
  assign pes_38_reset = reset;
  assign pes_38_io_cfg_en = cfgRegs_10[44]; // @[CGRA.scala 513:35]
  assign pes_38_io_cfg_addr = cfgRegs_10[43:32]; // @[CGRA.scala 514:35]
  assign pes_38_io_cfg_data = cfgRegs_10[31:0]; // @[CGRA.scala 515:35]
  assign pes_38_io_en = io_en_6; // @[CGRA.scala 377:27]
  assign pes_38_io_in_0 = gibs_42_io_ipinSE_0; // @[CGRA.scala 380:14]
  assign pes_38_io_in_1 = gibs_43_io_ipinSW_0; // @[CGRA.scala 384:14]
  assign pes_38_io_in_2 = gibs_51_io_ipinNE_0; // @[CGRA.scala 388:14]
  assign pes_38_io_in_3 = gibs_52_io_ipinNW_0; // @[CGRA.scala 392:14]
  assign pes_38_io_in_4 = gibs_42_io_ipinSE_1; // @[CGRA.scala 380:14]
  assign pes_38_io_in_5 = gibs_43_io_ipinSW_1; // @[CGRA.scala 384:14]
  assign pes_38_io_in_6 = gibs_51_io_ipinNE_1; // @[CGRA.scala 388:14]
  assign pes_38_io_in_7 = gibs_52_io_ipinNW_1; // @[CGRA.scala 392:14]
  assign pes_39_clock = clock;
  assign pes_39_reset = reset;
  assign pes_39_io_cfg_en = cfgRegs_10[44]; // @[CGRA.scala 513:35]
  assign pes_39_io_cfg_addr = cfgRegs_10[43:32]; // @[CGRA.scala 514:35]
  assign pes_39_io_cfg_data = cfgRegs_10[31:0]; // @[CGRA.scala 515:35]
  assign pes_39_io_en = io_en_7; // @[CGRA.scala 377:27]
  assign pes_39_io_in_0 = gibs_43_io_ipinSE_0; // @[CGRA.scala 380:14]
  assign pes_39_io_in_1 = gibs_44_io_ipinSW_0; // @[CGRA.scala 384:14]
  assign pes_39_io_in_2 = gibs_52_io_ipinNE_0; // @[CGRA.scala 388:14]
  assign pes_39_io_in_3 = gibs_53_io_ipinNW_0; // @[CGRA.scala 392:14]
  assign pes_39_io_in_4 = gibs_43_io_ipinSE_1; // @[CGRA.scala 380:14]
  assign pes_39_io_in_5 = gibs_44_io_ipinSW_1; // @[CGRA.scala 384:14]
  assign pes_39_io_in_6 = gibs_52_io_ipinNE_1; // @[CGRA.scala 388:14]
  assign pes_39_io_in_7 = gibs_53_io_ipinNW_1; // @[CGRA.scala 392:14]
  assign pes_40_clock = clock;
  assign pes_40_reset = reset;
  assign pes_40_io_cfg_en = cfgRegs_12[44]; // @[CGRA.scala 513:35]
  assign pes_40_io_cfg_addr = cfgRegs_12[43:32]; // @[CGRA.scala 514:35]
  assign pes_40_io_cfg_data = cfgRegs_12[31:0]; // @[CGRA.scala 515:35]
  assign pes_40_io_en = io_en_0; // @[CGRA.scala 377:27]
  assign pes_40_io_in_0 = gibs_45_io_ipinSE_0; // @[CGRA.scala 380:14]
  assign pes_40_io_in_1 = gibs_46_io_ipinSW_0; // @[CGRA.scala 384:14]
  assign pes_40_io_in_2 = gibs_54_io_ipinNE_0; // @[CGRA.scala 388:14]
  assign pes_40_io_in_3 = gibs_55_io_ipinNW_0; // @[CGRA.scala 392:14]
  assign pes_40_io_in_4 = gibs_45_io_ipinSE_1; // @[CGRA.scala 380:14]
  assign pes_40_io_in_5 = gibs_46_io_ipinSW_1; // @[CGRA.scala 384:14]
  assign pes_40_io_in_6 = gibs_54_io_ipinNE_1; // @[CGRA.scala 388:14]
  assign pes_40_io_in_7 = gibs_55_io_ipinNW_1; // @[CGRA.scala 392:14]
  assign pes_41_clock = clock;
  assign pes_41_reset = reset;
  assign pes_41_io_cfg_en = cfgRegs_12[44]; // @[CGRA.scala 513:35]
  assign pes_41_io_cfg_addr = cfgRegs_12[43:32]; // @[CGRA.scala 514:35]
  assign pes_41_io_cfg_data = cfgRegs_12[31:0]; // @[CGRA.scala 515:35]
  assign pes_41_io_en = io_en_1; // @[CGRA.scala 377:27]
  assign pes_41_io_in_0 = gibs_46_io_ipinSE_0; // @[CGRA.scala 380:14]
  assign pes_41_io_in_1 = gibs_47_io_ipinSW_0; // @[CGRA.scala 384:14]
  assign pes_41_io_in_2 = gibs_55_io_ipinNE_0; // @[CGRA.scala 388:14]
  assign pes_41_io_in_3 = gibs_56_io_ipinNW_0; // @[CGRA.scala 392:14]
  assign pes_41_io_in_4 = gibs_46_io_ipinSE_1; // @[CGRA.scala 380:14]
  assign pes_41_io_in_5 = gibs_47_io_ipinSW_1; // @[CGRA.scala 384:14]
  assign pes_41_io_in_6 = gibs_55_io_ipinNE_1; // @[CGRA.scala 388:14]
  assign pes_41_io_in_7 = gibs_56_io_ipinNW_1; // @[CGRA.scala 392:14]
  assign pes_42_clock = clock;
  assign pes_42_reset = reset;
  assign pes_42_io_cfg_en = cfgRegs_12[44]; // @[CGRA.scala 513:35]
  assign pes_42_io_cfg_addr = cfgRegs_12[43:32]; // @[CGRA.scala 514:35]
  assign pes_42_io_cfg_data = cfgRegs_12[31:0]; // @[CGRA.scala 515:35]
  assign pes_42_io_en = io_en_2; // @[CGRA.scala 377:27]
  assign pes_42_io_in_0 = gibs_47_io_ipinSE_0; // @[CGRA.scala 380:14]
  assign pes_42_io_in_1 = gibs_48_io_ipinSW_0; // @[CGRA.scala 384:14]
  assign pes_42_io_in_2 = gibs_56_io_ipinNE_0; // @[CGRA.scala 388:14]
  assign pes_42_io_in_3 = gibs_57_io_ipinNW_0; // @[CGRA.scala 392:14]
  assign pes_42_io_in_4 = gibs_47_io_ipinSE_1; // @[CGRA.scala 380:14]
  assign pes_42_io_in_5 = gibs_48_io_ipinSW_1; // @[CGRA.scala 384:14]
  assign pes_42_io_in_6 = gibs_56_io_ipinNE_1; // @[CGRA.scala 388:14]
  assign pes_42_io_in_7 = gibs_57_io_ipinNW_1; // @[CGRA.scala 392:14]
  assign pes_43_clock = clock;
  assign pes_43_reset = reset;
  assign pes_43_io_cfg_en = cfgRegs_12[44]; // @[CGRA.scala 513:35]
  assign pes_43_io_cfg_addr = cfgRegs_12[43:32]; // @[CGRA.scala 514:35]
  assign pes_43_io_cfg_data = cfgRegs_12[31:0]; // @[CGRA.scala 515:35]
  assign pes_43_io_en = io_en_3; // @[CGRA.scala 377:27]
  assign pes_43_io_in_0 = gibs_48_io_ipinSE_0; // @[CGRA.scala 380:14]
  assign pes_43_io_in_1 = gibs_49_io_ipinSW_0; // @[CGRA.scala 384:14]
  assign pes_43_io_in_2 = gibs_57_io_ipinNE_0; // @[CGRA.scala 388:14]
  assign pes_43_io_in_3 = gibs_58_io_ipinNW_0; // @[CGRA.scala 392:14]
  assign pes_43_io_in_4 = gibs_48_io_ipinSE_1; // @[CGRA.scala 380:14]
  assign pes_43_io_in_5 = gibs_49_io_ipinSW_1; // @[CGRA.scala 384:14]
  assign pes_43_io_in_6 = gibs_57_io_ipinNE_1; // @[CGRA.scala 388:14]
  assign pes_43_io_in_7 = gibs_58_io_ipinNW_1; // @[CGRA.scala 392:14]
  assign pes_44_clock = clock;
  assign pes_44_reset = reset;
  assign pes_44_io_cfg_en = cfgRegs_12[44]; // @[CGRA.scala 513:35]
  assign pes_44_io_cfg_addr = cfgRegs_12[43:32]; // @[CGRA.scala 514:35]
  assign pes_44_io_cfg_data = cfgRegs_12[31:0]; // @[CGRA.scala 515:35]
  assign pes_44_io_en = io_en_4; // @[CGRA.scala 377:27]
  assign pes_44_io_in_0 = gibs_49_io_ipinSE_0; // @[CGRA.scala 380:14]
  assign pes_44_io_in_1 = gibs_50_io_ipinSW_0; // @[CGRA.scala 384:14]
  assign pes_44_io_in_2 = gibs_58_io_ipinNE_0; // @[CGRA.scala 388:14]
  assign pes_44_io_in_3 = gibs_59_io_ipinNW_0; // @[CGRA.scala 392:14]
  assign pes_44_io_in_4 = gibs_49_io_ipinSE_1; // @[CGRA.scala 380:14]
  assign pes_44_io_in_5 = gibs_50_io_ipinSW_1; // @[CGRA.scala 384:14]
  assign pes_44_io_in_6 = gibs_58_io_ipinNE_1; // @[CGRA.scala 388:14]
  assign pes_44_io_in_7 = gibs_59_io_ipinNW_1; // @[CGRA.scala 392:14]
  assign pes_45_clock = clock;
  assign pes_45_reset = reset;
  assign pes_45_io_cfg_en = cfgRegs_12[44]; // @[CGRA.scala 513:35]
  assign pes_45_io_cfg_addr = cfgRegs_12[43:32]; // @[CGRA.scala 514:35]
  assign pes_45_io_cfg_data = cfgRegs_12[31:0]; // @[CGRA.scala 515:35]
  assign pes_45_io_en = io_en_5; // @[CGRA.scala 377:27]
  assign pes_45_io_in_0 = gibs_50_io_ipinSE_0; // @[CGRA.scala 380:14]
  assign pes_45_io_in_1 = gibs_51_io_ipinSW_0; // @[CGRA.scala 384:14]
  assign pes_45_io_in_2 = gibs_59_io_ipinNE_0; // @[CGRA.scala 388:14]
  assign pes_45_io_in_3 = gibs_60_io_ipinNW_0; // @[CGRA.scala 392:14]
  assign pes_45_io_in_4 = gibs_50_io_ipinSE_1; // @[CGRA.scala 380:14]
  assign pes_45_io_in_5 = gibs_51_io_ipinSW_1; // @[CGRA.scala 384:14]
  assign pes_45_io_in_6 = gibs_59_io_ipinNE_1; // @[CGRA.scala 388:14]
  assign pes_45_io_in_7 = gibs_60_io_ipinNW_1; // @[CGRA.scala 392:14]
  assign pes_46_clock = clock;
  assign pes_46_reset = reset;
  assign pes_46_io_cfg_en = cfgRegs_12[44]; // @[CGRA.scala 513:35]
  assign pes_46_io_cfg_addr = cfgRegs_12[43:32]; // @[CGRA.scala 514:35]
  assign pes_46_io_cfg_data = cfgRegs_12[31:0]; // @[CGRA.scala 515:35]
  assign pes_46_io_en = io_en_6; // @[CGRA.scala 377:27]
  assign pes_46_io_in_0 = gibs_51_io_ipinSE_0; // @[CGRA.scala 380:14]
  assign pes_46_io_in_1 = gibs_52_io_ipinSW_0; // @[CGRA.scala 384:14]
  assign pes_46_io_in_2 = gibs_60_io_ipinNE_0; // @[CGRA.scala 388:14]
  assign pes_46_io_in_3 = gibs_61_io_ipinNW_0; // @[CGRA.scala 392:14]
  assign pes_46_io_in_4 = gibs_51_io_ipinSE_1; // @[CGRA.scala 380:14]
  assign pes_46_io_in_5 = gibs_52_io_ipinSW_1; // @[CGRA.scala 384:14]
  assign pes_46_io_in_6 = gibs_60_io_ipinNE_1; // @[CGRA.scala 388:14]
  assign pes_46_io_in_7 = gibs_61_io_ipinNW_1; // @[CGRA.scala 392:14]
  assign pes_47_clock = clock;
  assign pes_47_reset = reset;
  assign pes_47_io_cfg_en = cfgRegs_12[44]; // @[CGRA.scala 513:35]
  assign pes_47_io_cfg_addr = cfgRegs_12[43:32]; // @[CGRA.scala 514:35]
  assign pes_47_io_cfg_data = cfgRegs_12[31:0]; // @[CGRA.scala 515:35]
  assign pes_47_io_en = io_en_7; // @[CGRA.scala 377:27]
  assign pes_47_io_in_0 = gibs_52_io_ipinSE_0; // @[CGRA.scala 380:14]
  assign pes_47_io_in_1 = gibs_53_io_ipinSW_0; // @[CGRA.scala 384:14]
  assign pes_47_io_in_2 = gibs_61_io_ipinNE_0; // @[CGRA.scala 388:14]
  assign pes_47_io_in_3 = gibs_62_io_ipinNW_0; // @[CGRA.scala 392:14]
  assign pes_47_io_in_4 = gibs_52_io_ipinSE_1; // @[CGRA.scala 380:14]
  assign pes_47_io_in_5 = gibs_53_io_ipinSW_1; // @[CGRA.scala 384:14]
  assign pes_47_io_in_6 = gibs_61_io_ipinNE_1; // @[CGRA.scala 388:14]
  assign pes_47_io_in_7 = gibs_62_io_ipinNW_1; // @[CGRA.scala 392:14]
  assign pes_48_clock = clock;
  assign pes_48_reset = reset;
  assign pes_48_io_cfg_en = cfgRegs_14[44]; // @[CGRA.scala 513:35]
  assign pes_48_io_cfg_addr = cfgRegs_14[43:32]; // @[CGRA.scala 514:35]
  assign pes_48_io_cfg_data = cfgRegs_14[31:0]; // @[CGRA.scala 515:35]
  assign pes_48_io_en = io_en_0; // @[CGRA.scala 377:27]
  assign pes_48_io_in_0 = gibs_54_io_ipinSE_0; // @[CGRA.scala 380:14]
  assign pes_48_io_in_1 = gibs_55_io_ipinSW_0; // @[CGRA.scala 384:14]
  assign pes_48_io_in_2 = gibs_63_io_ipinNE_0; // @[CGRA.scala 388:14]
  assign pes_48_io_in_3 = gibs_64_io_ipinNW_0; // @[CGRA.scala 392:14]
  assign pes_48_io_in_4 = gibs_54_io_ipinSE_1; // @[CGRA.scala 380:14]
  assign pes_48_io_in_5 = gibs_55_io_ipinSW_1; // @[CGRA.scala 384:14]
  assign pes_48_io_in_6 = gibs_63_io_ipinNE_1; // @[CGRA.scala 388:14]
  assign pes_48_io_in_7 = gibs_64_io_ipinNW_1; // @[CGRA.scala 392:14]
  assign pes_49_clock = clock;
  assign pes_49_reset = reset;
  assign pes_49_io_cfg_en = cfgRegs_14[44]; // @[CGRA.scala 513:35]
  assign pes_49_io_cfg_addr = cfgRegs_14[43:32]; // @[CGRA.scala 514:35]
  assign pes_49_io_cfg_data = cfgRegs_14[31:0]; // @[CGRA.scala 515:35]
  assign pes_49_io_en = io_en_1; // @[CGRA.scala 377:27]
  assign pes_49_io_in_0 = gibs_55_io_ipinSE_0; // @[CGRA.scala 380:14]
  assign pes_49_io_in_1 = gibs_56_io_ipinSW_0; // @[CGRA.scala 384:14]
  assign pes_49_io_in_2 = gibs_64_io_ipinNE_0; // @[CGRA.scala 388:14]
  assign pes_49_io_in_3 = gibs_65_io_ipinNW_0; // @[CGRA.scala 392:14]
  assign pes_49_io_in_4 = gibs_55_io_ipinSE_1; // @[CGRA.scala 380:14]
  assign pes_49_io_in_5 = gibs_56_io_ipinSW_1; // @[CGRA.scala 384:14]
  assign pes_49_io_in_6 = gibs_64_io_ipinNE_1; // @[CGRA.scala 388:14]
  assign pes_49_io_in_7 = gibs_65_io_ipinNW_1; // @[CGRA.scala 392:14]
  assign pes_50_clock = clock;
  assign pes_50_reset = reset;
  assign pes_50_io_cfg_en = cfgRegs_14[44]; // @[CGRA.scala 513:35]
  assign pes_50_io_cfg_addr = cfgRegs_14[43:32]; // @[CGRA.scala 514:35]
  assign pes_50_io_cfg_data = cfgRegs_14[31:0]; // @[CGRA.scala 515:35]
  assign pes_50_io_en = io_en_2; // @[CGRA.scala 377:27]
  assign pes_50_io_in_0 = gibs_56_io_ipinSE_0; // @[CGRA.scala 380:14]
  assign pes_50_io_in_1 = gibs_57_io_ipinSW_0; // @[CGRA.scala 384:14]
  assign pes_50_io_in_2 = gibs_65_io_ipinNE_0; // @[CGRA.scala 388:14]
  assign pes_50_io_in_3 = gibs_66_io_ipinNW_0; // @[CGRA.scala 392:14]
  assign pes_50_io_in_4 = gibs_56_io_ipinSE_1; // @[CGRA.scala 380:14]
  assign pes_50_io_in_5 = gibs_57_io_ipinSW_1; // @[CGRA.scala 384:14]
  assign pes_50_io_in_6 = gibs_65_io_ipinNE_1; // @[CGRA.scala 388:14]
  assign pes_50_io_in_7 = gibs_66_io_ipinNW_1; // @[CGRA.scala 392:14]
  assign pes_51_clock = clock;
  assign pes_51_reset = reset;
  assign pes_51_io_cfg_en = cfgRegs_14[44]; // @[CGRA.scala 513:35]
  assign pes_51_io_cfg_addr = cfgRegs_14[43:32]; // @[CGRA.scala 514:35]
  assign pes_51_io_cfg_data = cfgRegs_14[31:0]; // @[CGRA.scala 515:35]
  assign pes_51_io_en = io_en_3; // @[CGRA.scala 377:27]
  assign pes_51_io_in_0 = gibs_57_io_ipinSE_0; // @[CGRA.scala 380:14]
  assign pes_51_io_in_1 = gibs_58_io_ipinSW_0; // @[CGRA.scala 384:14]
  assign pes_51_io_in_2 = gibs_66_io_ipinNE_0; // @[CGRA.scala 388:14]
  assign pes_51_io_in_3 = gibs_67_io_ipinNW_0; // @[CGRA.scala 392:14]
  assign pes_51_io_in_4 = gibs_57_io_ipinSE_1; // @[CGRA.scala 380:14]
  assign pes_51_io_in_5 = gibs_58_io_ipinSW_1; // @[CGRA.scala 384:14]
  assign pes_51_io_in_6 = gibs_66_io_ipinNE_1; // @[CGRA.scala 388:14]
  assign pes_51_io_in_7 = gibs_67_io_ipinNW_1; // @[CGRA.scala 392:14]
  assign pes_52_clock = clock;
  assign pes_52_reset = reset;
  assign pes_52_io_cfg_en = cfgRegs_14[44]; // @[CGRA.scala 513:35]
  assign pes_52_io_cfg_addr = cfgRegs_14[43:32]; // @[CGRA.scala 514:35]
  assign pes_52_io_cfg_data = cfgRegs_14[31:0]; // @[CGRA.scala 515:35]
  assign pes_52_io_en = io_en_4; // @[CGRA.scala 377:27]
  assign pes_52_io_in_0 = gibs_58_io_ipinSE_0; // @[CGRA.scala 380:14]
  assign pes_52_io_in_1 = gibs_59_io_ipinSW_0; // @[CGRA.scala 384:14]
  assign pes_52_io_in_2 = gibs_67_io_ipinNE_0; // @[CGRA.scala 388:14]
  assign pes_52_io_in_3 = gibs_68_io_ipinNW_0; // @[CGRA.scala 392:14]
  assign pes_52_io_in_4 = gibs_58_io_ipinSE_1; // @[CGRA.scala 380:14]
  assign pes_52_io_in_5 = gibs_59_io_ipinSW_1; // @[CGRA.scala 384:14]
  assign pes_52_io_in_6 = gibs_67_io_ipinNE_1; // @[CGRA.scala 388:14]
  assign pes_52_io_in_7 = gibs_68_io_ipinNW_1; // @[CGRA.scala 392:14]
  assign pes_53_clock = clock;
  assign pes_53_reset = reset;
  assign pes_53_io_cfg_en = cfgRegs_14[44]; // @[CGRA.scala 513:35]
  assign pes_53_io_cfg_addr = cfgRegs_14[43:32]; // @[CGRA.scala 514:35]
  assign pes_53_io_cfg_data = cfgRegs_14[31:0]; // @[CGRA.scala 515:35]
  assign pes_53_io_en = io_en_5; // @[CGRA.scala 377:27]
  assign pes_53_io_in_0 = gibs_59_io_ipinSE_0; // @[CGRA.scala 380:14]
  assign pes_53_io_in_1 = gibs_60_io_ipinSW_0; // @[CGRA.scala 384:14]
  assign pes_53_io_in_2 = gibs_68_io_ipinNE_0; // @[CGRA.scala 388:14]
  assign pes_53_io_in_3 = gibs_69_io_ipinNW_0; // @[CGRA.scala 392:14]
  assign pes_53_io_in_4 = gibs_59_io_ipinSE_1; // @[CGRA.scala 380:14]
  assign pes_53_io_in_5 = gibs_60_io_ipinSW_1; // @[CGRA.scala 384:14]
  assign pes_53_io_in_6 = gibs_68_io_ipinNE_1; // @[CGRA.scala 388:14]
  assign pes_53_io_in_7 = gibs_69_io_ipinNW_1; // @[CGRA.scala 392:14]
  assign pes_54_clock = clock;
  assign pes_54_reset = reset;
  assign pes_54_io_cfg_en = cfgRegs_14[44]; // @[CGRA.scala 513:35]
  assign pes_54_io_cfg_addr = cfgRegs_14[43:32]; // @[CGRA.scala 514:35]
  assign pes_54_io_cfg_data = cfgRegs_14[31:0]; // @[CGRA.scala 515:35]
  assign pes_54_io_en = io_en_6; // @[CGRA.scala 377:27]
  assign pes_54_io_in_0 = gibs_60_io_ipinSE_0; // @[CGRA.scala 380:14]
  assign pes_54_io_in_1 = gibs_61_io_ipinSW_0; // @[CGRA.scala 384:14]
  assign pes_54_io_in_2 = gibs_69_io_ipinNE_0; // @[CGRA.scala 388:14]
  assign pes_54_io_in_3 = gibs_70_io_ipinNW_0; // @[CGRA.scala 392:14]
  assign pes_54_io_in_4 = gibs_60_io_ipinSE_1; // @[CGRA.scala 380:14]
  assign pes_54_io_in_5 = gibs_61_io_ipinSW_1; // @[CGRA.scala 384:14]
  assign pes_54_io_in_6 = gibs_69_io_ipinNE_1; // @[CGRA.scala 388:14]
  assign pes_54_io_in_7 = gibs_70_io_ipinNW_1; // @[CGRA.scala 392:14]
  assign pes_55_clock = clock;
  assign pes_55_reset = reset;
  assign pes_55_io_cfg_en = cfgRegs_14[44]; // @[CGRA.scala 513:35]
  assign pes_55_io_cfg_addr = cfgRegs_14[43:32]; // @[CGRA.scala 514:35]
  assign pes_55_io_cfg_data = cfgRegs_14[31:0]; // @[CGRA.scala 515:35]
  assign pes_55_io_en = io_en_7; // @[CGRA.scala 377:27]
  assign pes_55_io_in_0 = gibs_61_io_ipinSE_0; // @[CGRA.scala 380:14]
  assign pes_55_io_in_1 = gibs_62_io_ipinSW_0; // @[CGRA.scala 384:14]
  assign pes_55_io_in_2 = gibs_70_io_ipinNE_0; // @[CGRA.scala 388:14]
  assign pes_55_io_in_3 = gibs_71_io_ipinNW_0; // @[CGRA.scala 392:14]
  assign pes_55_io_in_4 = gibs_61_io_ipinSE_1; // @[CGRA.scala 380:14]
  assign pes_55_io_in_5 = gibs_62_io_ipinSW_1; // @[CGRA.scala 384:14]
  assign pes_55_io_in_6 = gibs_70_io_ipinNE_1; // @[CGRA.scala 388:14]
  assign pes_55_io_in_7 = gibs_71_io_ipinNW_1; // @[CGRA.scala 392:14]
  assign pes_56_clock = clock;
  assign pes_56_reset = reset;
  assign pes_56_io_cfg_en = cfgRegs_16[44]; // @[CGRA.scala 513:35]
  assign pes_56_io_cfg_addr = cfgRegs_16[43:32]; // @[CGRA.scala 514:35]
  assign pes_56_io_cfg_data = cfgRegs_16[31:0]; // @[CGRA.scala 515:35]
  assign pes_56_io_en = io_en_0; // @[CGRA.scala 377:27]
  assign pes_56_io_in_0 = gibs_63_io_ipinSE_0; // @[CGRA.scala 380:14]
  assign pes_56_io_in_1 = gibs_64_io_ipinSW_0; // @[CGRA.scala 384:14]
  assign pes_56_io_in_2 = gibs_72_io_ipinNE_0; // @[CGRA.scala 388:14]
  assign pes_56_io_in_3 = gibs_73_io_ipinNW_0; // @[CGRA.scala 392:14]
  assign pes_56_io_in_4 = gibs_63_io_ipinSE_1; // @[CGRA.scala 380:14]
  assign pes_56_io_in_5 = gibs_64_io_ipinSW_1; // @[CGRA.scala 384:14]
  assign pes_56_io_in_6 = gibs_72_io_ipinNE_1; // @[CGRA.scala 388:14]
  assign pes_56_io_in_7 = gibs_73_io_ipinNW_1; // @[CGRA.scala 392:14]
  assign pes_57_clock = clock;
  assign pes_57_reset = reset;
  assign pes_57_io_cfg_en = cfgRegs_16[44]; // @[CGRA.scala 513:35]
  assign pes_57_io_cfg_addr = cfgRegs_16[43:32]; // @[CGRA.scala 514:35]
  assign pes_57_io_cfg_data = cfgRegs_16[31:0]; // @[CGRA.scala 515:35]
  assign pes_57_io_en = io_en_1; // @[CGRA.scala 377:27]
  assign pes_57_io_in_0 = gibs_64_io_ipinSE_0; // @[CGRA.scala 380:14]
  assign pes_57_io_in_1 = gibs_65_io_ipinSW_0; // @[CGRA.scala 384:14]
  assign pes_57_io_in_2 = gibs_73_io_ipinNE_0; // @[CGRA.scala 388:14]
  assign pes_57_io_in_3 = gibs_74_io_ipinNW_0; // @[CGRA.scala 392:14]
  assign pes_57_io_in_4 = gibs_64_io_ipinSE_1; // @[CGRA.scala 380:14]
  assign pes_57_io_in_5 = gibs_65_io_ipinSW_1; // @[CGRA.scala 384:14]
  assign pes_57_io_in_6 = gibs_73_io_ipinNE_1; // @[CGRA.scala 388:14]
  assign pes_57_io_in_7 = gibs_74_io_ipinNW_1; // @[CGRA.scala 392:14]
  assign pes_58_clock = clock;
  assign pes_58_reset = reset;
  assign pes_58_io_cfg_en = cfgRegs_16[44]; // @[CGRA.scala 513:35]
  assign pes_58_io_cfg_addr = cfgRegs_16[43:32]; // @[CGRA.scala 514:35]
  assign pes_58_io_cfg_data = cfgRegs_16[31:0]; // @[CGRA.scala 515:35]
  assign pes_58_io_en = io_en_2; // @[CGRA.scala 377:27]
  assign pes_58_io_in_0 = gibs_65_io_ipinSE_0; // @[CGRA.scala 380:14]
  assign pes_58_io_in_1 = gibs_66_io_ipinSW_0; // @[CGRA.scala 384:14]
  assign pes_58_io_in_2 = gibs_74_io_ipinNE_0; // @[CGRA.scala 388:14]
  assign pes_58_io_in_3 = gibs_75_io_ipinNW_0; // @[CGRA.scala 392:14]
  assign pes_58_io_in_4 = gibs_65_io_ipinSE_1; // @[CGRA.scala 380:14]
  assign pes_58_io_in_5 = gibs_66_io_ipinSW_1; // @[CGRA.scala 384:14]
  assign pes_58_io_in_6 = gibs_74_io_ipinNE_1; // @[CGRA.scala 388:14]
  assign pes_58_io_in_7 = gibs_75_io_ipinNW_1; // @[CGRA.scala 392:14]
  assign pes_59_clock = clock;
  assign pes_59_reset = reset;
  assign pes_59_io_cfg_en = cfgRegs_16[44]; // @[CGRA.scala 513:35]
  assign pes_59_io_cfg_addr = cfgRegs_16[43:32]; // @[CGRA.scala 514:35]
  assign pes_59_io_cfg_data = cfgRegs_16[31:0]; // @[CGRA.scala 515:35]
  assign pes_59_io_en = io_en_3; // @[CGRA.scala 377:27]
  assign pes_59_io_in_0 = gibs_66_io_ipinSE_0; // @[CGRA.scala 380:14]
  assign pes_59_io_in_1 = gibs_67_io_ipinSW_0; // @[CGRA.scala 384:14]
  assign pes_59_io_in_2 = gibs_75_io_ipinNE_0; // @[CGRA.scala 388:14]
  assign pes_59_io_in_3 = gibs_76_io_ipinNW_0; // @[CGRA.scala 392:14]
  assign pes_59_io_in_4 = gibs_66_io_ipinSE_1; // @[CGRA.scala 380:14]
  assign pes_59_io_in_5 = gibs_67_io_ipinSW_1; // @[CGRA.scala 384:14]
  assign pes_59_io_in_6 = gibs_75_io_ipinNE_1; // @[CGRA.scala 388:14]
  assign pes_59_io_in_7 = gibs_76_io_ipinNW_1; // @[CGRA.scala 392:14]
  assign pes_60_clock = clock;
  assign pes_60_reset = reset;
  assign pes_60_io_cfg_en = cfgRegs_16[44]; // @[CGRA.scala 513:35]
  assign pes_60_io_cfg_addr = cfgRegs_16[43:32]; // @[CGRA.scala 514:35]
  assign pes_60_io_cfg_data = cfgRegs_16[31:0]; // @[CGRA.scala 515:35]
  assign pes_60_io_en = io_en_4; // @[CGRA.scala 377:27]
  assign pes_60_io_in_0 = gibs_67_io_ipinSE_0; // @[CGRA.scala 380:14]
  assign pes_60_io_in_1 = gibs_68_io_ipinSW_0; // @[CGRA.scala 384:14]
  assign pes_60_io_in_2 = gibs_76_io_ipinNE_0; // @[CGRA.scala 388:14]
  assign pes_60_io_in_3 = gibs_77_io_ipinNW_0; // @[CGRA.scala 392:14]
  assign pes_60_io_in_4 = gibs_67_io_ipinSE_1; // @[CGRA.scala 380:14]
  assign pes_60_io_in_5 = gibs_68_io_ipinSW_1; // @[CGRA.scala 384:14]
  assign pes_60_io_in_6 = gibs_76_io_ipinNE_1; // @[CGRA.scala 388:14]
  assign pes_60_io_in_7 = gibs_77_io_ipinNW_1; // @[CGRA.scala 392:14]
  assign pes_61_clock = clock;
  assign pes_61_reset = reset;
  assign pes_61_io_cfg_en = cfgRegs_16[44]; // @[CGRA.scala 513:35]
  assign pes_61_io_cfg_addr = cfgRegs_16[43:32]; // @[CGRA.scala 514:35]
  assign pes_61_io_cfg_data = cfgRegs_16[31:0]; // @[CGRA.scala 515:35]
  assign pes_61_io_en = io_en_5; // @[CGRA.scala 377:27]
  assign pes_61_io_in_0 = gibs_68_io_ipinSE_0; // @[CGRA.scala 380:14]
  assign pes_61_io_in_1 = gibs_69_io_ipinSW_0; // @[CGRA.scala 384:14]
  assign pes_61_io_in_2 = gibs_77_io_ipinNE_0; // @[CGRA.scala 388:14]
  assign pes_61_io_in_3 = gibs_78_io_ipinNW_0; // @[CGRA.scala 392:14]
  assign pes_61_io_in_4 = gibs_68_io_ipinSE_1; // @[CGRA.scala 380:14]
  assign pes_61_io_in_5 = gibs_69_io_ipinSW_1; // @[CGRA.scala 384:14]
  assign pes_61_io_in_6 = gibs_77_io_ipinNE_1; // @[CGRA.scala 388:14]
  assign pes_61_io_in_7 = gibs_78_io_ipinNW_1; // @[CGRA.scala 392:14]
  assign pes_62_clock = clock;
  assign pes_62_reset = reset;
  assign pes_62_io_cfg_en = cfgRegs_16[44]; // @[CGRA.scala 513:35]
  assign pes_62_io_cfg_addr = cfgRegs_16[43:32]; // @[CGRA.scala 514:35]
  assign pes_62_io_cfg_data = cfgRegs_16[31:0]; // @[CGRA.scala 515:35]
  assign pes_62_io_en = io_en_6; // @[CGRA.scala 377:27]
  assign pes_62_io_in_0 = gibs_69_io_ipinSE_0; // @[CGRA.scala 380:14]
  assign pes_62_io_in_1 = gibs_70_io_ipinSW_0; // @[CGRA.scala 384:14]
  assign pes_62_io_in_2 = gibs_78_io_ipinNE_0; // @[CGRA.scala 388:14]
  assign pes_62_io_in_3 = gibs_79_io_ipinNW_0; // @[CGRA.scala 392:14]
  assign pes_62_io_in_4 = gibs_69_io_ipinSE_1; // @[CGRA.scala 380:14]
  assign pes_62_io_in_5 = gibs_70_io_ipinSW_1; // @[CGRA.scala 384:14]
  assign pes_62_io_in_6 = gibs_78_io_ipinNE_1; // @[CGRA.scala 388:14]
  assign pes_62_io_in_7 = gibs_79_io_ipinNW_1; // @[CGRA.scala 392:14]
  assign pes_63_clock = clock;
  assign pes_63_reset = reset;
  assign pes_63_io_cfg_en = cfgRegs_16[44]; // @[CGRA.scala 513:35]
  assign pes_63_io_cfg_addr = cfgRegs_16[43:32]; // @[CGRA.scala 514:35]
  assign pes_63_io_cfg_data = cfgRegs_16[31:0]; // @[CGRA.scala 515:35]
  assign pes_63_io_en = io_en_7; // @[CGRA.scala 377:27]
  assign pes_63_io_in_0 = gibs_70_io_ipinSE_0; // @[CGRA.scala 380:14]
  assign pes_63_io_in_1 = gibs_71_io_ipinSW_0; // @[CGRA.scala 384:14]
  assign pes_63_io_in_2 = gibs_79_io_ipinNE_0; // @[CGRA.scala 388:14]
  assign pes_63_io_in_3 = gibs_80_io_ipinNW_0; // @[CGRA.scala 392:14]
  assign pes_63_io_in_4 = gibs_70_io_ipinSE_1; // @[CGRA.scala 380:14]
  assign pes_63_io_in_5 = gibs_71_io_ipinSW_1; // @[CGRA.scala 384:14]
  assign pes_63_io_in_6 = gibs_79_io_ipinNE_1; // @[CGRA.scala 388:14]
  assign pes_63_io_in_7 = gibs_80_io_ipinNW_1; // @[CGRA.scala 392:14]
  assign gibs_0_clock = clock;
  assign gibs_0_reset = reset;
  assign gibs_0_io_cfg_en = cfgRegs_1[44]; // @[CGRA.scala 509:38]
  assign gibs_0_io_cfg_addr = cfgRegs_1[43:32]; // @[CGRA.scala 510:38]
  assign gibs_0_io_cfg_data = cfgRegs_1[31:0]; // @[CGRA.scala 511:38]
  assign gibs_0_io_opinNE_0 = ibs_0_io_out_0; // @[CGRA.scala 326:35]
  assign gibs_0_io_opinSE_0 = pes_0_io_out_0; // @[CGRA.scala 398:41]
  assign gibs_0_io_itrackE_0 = gibs_1_io_otrackW_0; // @[CGRA.scala 451:16]
  assign gibs_0_io_itrackS_0 = gibs_9_io_otrackN_0; // @[CGRA.scala 421:16]
  assign gibs_1_clock = clock;
  assign gibs_1_reset = reset;
  assign gibs_1_io_cfg_en = cfgRegs_1[44]; // @[CGRA.scala 509:38]
  assign gibs_1_io_cfg_addr = cfgRegs_1[43:32]; // @[CGRA.scala 510:38]
  assign gibs_1_io_cfg_data = cfgRegs_1[31:0]; // @[CGRA.scala 511:38]
  assign gibs_1_io_opinNW_0 = ibs_0_io_out_0; // @[CGRA.scala 327:37]
  assign gibs_1_io_opinNE_0 = ibs_1_io_out_0; // @[CGRA.scala 326:35]
  assign gibs_1_io_opinSE_0 = pes_1_io_out_0; // @[CGRA.scala 398:41]
  assign gibs_1_io_opinSW_0 = pes_0_io_out_0; // @[CGRA.scala 399:43]
  assign gibs_1_io_itrackW_0 = gibs_0_io_otrackE_0; // @[CGRA.scala 466:16]
  assign gibs_1_io_itrackE_0 = gibs_2_io_otrackW_0; // @[CGRA.scala 472:16]
  assign gibs_1_io_itrackS_0 = gibs_10_io_otrackN_0; // @[CGRA.scala 421:16]
  assign gibs_2_clock = clock;
  assign gibs_2_reset = reset;
  assign gibs_2_io_cfg_en = cfgRegs_1[44]; // @[CGRA.scala 509:38]
  assign gibs_2_io_cfg_addr = cfgRegs_1[43:32]; // @[CGRA.scala 510:38]
  assign gibs_2_io_cfg_data = cfgRegs_1[31:0]; // @[CGRA.scala 511:38]
  assign gibs_2_io_opinNW_0 = ibs_1_io_out_0; // @[CGRA.scala 327:37]
  assign gibs_2_io_opinNE_0 = ibs_2_io_out_0; // @[CGRA.scala 326:35]
  assign gibs_2_io_opinSE_0 = pes_2_io_out_0; // @[CGRA.scala 398:41]
  assign gibs_2_io_opinSW_0 = pes_1_io_out_0; // @[CGRA.scala 399:43]
  assign gibs_2_io_itrackW_0 = gibs_1_io_otrackE_0; // @[CGRA.scala 466:16]
  assign gibs_2_io_itrackE_0 = gibs_3_io_otrackW_0; // @[CGRA.scala 472:16]
  assign gibs_2_io_itrackS_0 = gibs_11_io_otrackN_0; // @[CGRA.scala 421:16]
  assign gibs_3_clock = clock;
  assign gibs_3_reset = reset;
  assign gibs_3_io_cfg_en = cfgRegs_1[44]; // @[CGRA.scala 509:38]
  assign gibs_3_io_cfg_addr = cfgRegs_1[43:32]; // @[CGRA.scala 510:38]
  assign gibs_3_io_cfg_data = cfgRegs_1[31:0]; // @[CGRA.scala 511:38]
  assign gibs_3_io_opinNW_0 = ibs_2_io_out_0; // @[CGRA.scala 327:37]
  assign gibs_3_io_opinNE_0 = ibs_3_io_out_0; // @[CGRA.scala 326:35]
  assign gibs_3_io_opinSE_0 = pes_3_io_out_0; // @[CGRA.scala 398:41]
  assign gibs_3_io_opinSW_0 = pes_2_io_out_0; // @[CGRA.scala 399:43]
  assign gibs_3_io_itrackW_0 = gibs_2_io_otrackE_0; // @[CGRA.scala 466:16]
  assign gibs_3_io_itrackE_0 = gibs_4_io_otrackW_0; // @[CGRA.scala 472:16]
  assign gibs_3_io_itrackS_0 = gibs_12_io_otrackN_0; // @[CGRA.scala 421:16]
  assign gibs_4_clock = clock;
  assign gibs_4_reset = reset;
  assign gibs_4_io_cfg_en = cfgRegs_1[44]; // @[CGRA.scala 509:38]
  assign gibs_4_io_cfg_addr = cfgRegs_1[43:32]; // @[CGRA.scala 510:38]
  assign gibs_4_io_cfg_data = cfgRegs_1[31:0]; // @[CGRA.scala 511:38]
  assign gibs_4_io_opinNW_0 = ibs_3_io_out_0; // @[CGRA.scala 327:37]
  assign gibs_4_io_opinNE_0 = ibs_4_io_out_0; // @[CGRA.scala 326:35]
  assign gibs_4_io_opinSE_0 = pes_4_io_out_0; // @[CGRA.scala 398:41]
  assign gibs_4_io_opinSW_0 = pes_3_io_out_0; // @[CGRA.scala 399:43]
  assign gibs_4_io_itrackW_0 = gibs_3_io_otrackE_0; // @[CGRA.scala 466:16]
  assign gibs_4_io_itrackE_0 = gibs_5_io_otrackW_0; // @[CGRA.scala 472:16]
  assign gibs_4_io_itrackS_0 = gibs_13_io_otrackN_0; // @[CGRA.scala 421:16]
  assign gibs_5_clock = clock;
  assign gibs_5_reset = reset;
  assign gibs_5_io_cfg_en = cfgRegs_1[44]; // @[CGRA.scala 509:38]
  assign gibs_5_io_cfg_addr = cfgRegs_1[43:32]; // @[CGRA.scala 510:38]
  assign gibs_5_io_cfg_data = cfgRegs_1[31:0]; // @[CGRA.scala 511:38]
  assign gibs_5_io_opinNW_0 = ibs_4_io_out_0; // @[CGRA.scala 327:37]
  assign gibs_5_io_opinNE_0 = ibs_5_io_out_0; // @[CGRA.scala 326:35]
  assign gibs_5_io_opinSE_0 = pes_5_io_out_0; // @[CGRA.scala 398:41]
  assign gibs_5_io_opinSW_0 = pes_4_io_out_0; // @[CGRA.scala 399:43]
  assign gibs_5_io_itrackW_0 = gibs_4_io_otrackE_0; // @[CGRA.scala 466:16]
  assign gibs_5_io_itrackE_0 = gibs_6_io_otrackW_0; // @[CGRA.scala 472:16]
  assign gibs_5_io_itrackS_0 = gibs_14_io_otrackN_0; // @[CGRA.scala 421:16]
  assign gibs_6_clock = clock;
  assign gibs_6_reset = reset;
  assign gibs_6_io_cfg_en = cfgRegs_1[44]; // @[CGRA.scala 509:38]
  assign gibs_6_io_cfg_addr = cfgRegs_1[43:32]; // @[CGRA.scala 510:38]
  assign gibs_6_io_cfg_data = cfgRegs_1[31:0]; // @[CGRA.scala 511:38]
  assign gibs_6_io_opinNW_0 = ibs_5_io_out_0; // @[CGRA.scala 327:37]
  assign gibs_6_io_opinNE_0 = ibs_6_io_out_0; // @[CGRA.scala 326:35]
  assign gibs_6_io_opinSE_0 = pes_6_io_out_0; // @[CGRA.scala 398:41]
  assign gibs_6_io_opinSW_0 = pes_5_io_out_0; // @[CGRA.scala 399:43]
  assign gibs_6_io_itrackW_0 = gibs_5_io_otrackE_0; // @[CGRA.scala 466:16]
  assign gibs_6_io_itrackE_0 = gibs_7_io_otrackW_0; // @[CGRA.scala 472:16]
  assign gibs_6_io_itrackS_0 = gibs_15_io_otrackN_0; // @[CGRA.scala 421:16]
  assign gibs_7_clock = clock;
  assign gibs_7_reset = reset;
  assign gibs_7_io_cfg_en = cfgRegs_1[44]; // @[CGRA.scala 509:38]
  assign gibs_7_io_cfg_addr = cfgRegs_1[43:32]; // @[CGRA.scala 510:38]
  assign gibs_7_io_cfg_data = cfgRegs_1[31:0]; // @[CGRA.scala 511:38]
  assign gibs_7_io_opinNW_0 = ibs_6_io_out_0; // @[CGRA.scala 327:37]
  assign gibs_7_io_opinNE_0 = ibs_7_io_out_0; // @[CGRA.scala 326:35]
  assign gibs_7_io_opinSE_0 = pes_7_io_out_0; // @[CGRA.scala 398:41]
  assign gibs_7_io_opinSW_0 = pes_6_io_out_0; // @[CGRA.scala 399:43]
  assign gibs_7_io_itrackW_0 = gibs_6_io_otrackE_0; // @[CGRA.scala 466:16]
  assign gibs_7_io_itrackE_0 = gibs_8_io_otrackW_0; // @[CGRA.scala 472:16]
  assign gibs_7_io_itrackS_0 = gibs_16_io_otrackN_0; // @[CGRA.scala 421:16]
  assign gibs_8_clock = clock;
  assign gibs_8_reset = reset;
  assign gibs_8_io_cfg_en = cfgRegs_1[44]; // @[CGRA.scala 509:38]
  assign gibs_8_io_cfg_addr = cfgRegs_1[43:32]; // @[CGRA.scala 510:38]
  assign gibs_8_io_cfg_data = cfgRegs_1[31:0]; // @[CGRA.scala 511:38]
  assign gibs_8_io_opinNW_0 = ibs_7_io_out_0; // @[CGRA.scala 327:37]
  assign gibs_8_io_opinSW_0 = pes_7_io_out_0; // @[CGRA.scala 399:43]
  assign gibs_8_io_itrackW_0 = gibs_7_io_otrackE_0; // @[CGRA.scala 459:16]
  assign gibs_8_io_itrackS_0 = gibs_17_io_otrackN_0; // @[CGRA.scala 421:16]
  assign gibs_9_clock = clock;
  assign gibs_9_reset = reset;
  assign gibs_9_io_cfg_en = cfgRegs_3[44]; // @[CGRA.scala 509:38]
  assign gibs_9_io_cfg_addr = cfgRegs_3[43:32]; // @[CGRA.scala 510:38]
  assign gibs_9_io_cfg_data = cfgRegs_3[31:0]; // @[CGRA.scala 511:38]
  assign gibs_9_io_opinNE_0 = pes_0_io_out_0; // @[CGRA.scala 400:45]
  assign gibs_9_io_opinSE_0 = pes_8_io_out_0; // @[CGRA.scala 398:41]
  assign gibs_9_io_itrackN_0 = gibs_0_io_otrackS_0; // @[CGRA.scala 436:16]
  assign gibs_9_io_itrackE_0 = gibs_10_io_otrackW_0; // @[CGRA.scala 451:16]
  assign gibs_9_io_itrackS_0 = gibs_18_io_otrackN_0; // @[CGRA.scala 442:16]
  assign gibs_10_clock = clock;
  assign gibs_10_reset = reset;
  assign gibs_10_io_cfg_en = cfgRegs_3[44]; // @[CGRA.scala 509:38]
  assign gibs_10_io_cfg_addr = cfgRegs_3[43:32]; // @[CGRA.scala 510:38]
  assign gibs_10_io_cfg_data = cfgRegs_3[31:0]; // @[CGRA.scala 511:38]
  assign gibs_10_io_opinNW_0 = pes_0_io_out_0; // @[CGRA.scala 401:47]
  assign gibs_10_io_opinNE_0 = pes_1_io_out_0; // @[CGRA.scala 400:45]
  assign gibs_10_io_opinSE_0 = pes_9_io_out_0; // @[CGRA.scala 398:41]
  assign gibs_10_io_opinSW_0 = pes_8_io_out_0; // @[CGRA.scala 399:43]
  assign gibs_10_io_itrackW_0 = gibs_9_io_otrackE_0; // @[CGRA.scala 466:16]
  assign gibs_10_io_itrackN_0 = gibs_1_io_otrackS_0; // @[CGRA.scala 436:16]
  assign gibs_10_io_itrackE_0 = gibs_11_io_otrackW_0; // @[CGRA.scala 472:16]
  assign gibs_10_io_itrackS_0 = gibs_19_io_otrackN_0; // @[CGRA.scala 442:16]
  assign gibs_11_clock = clock;
  assign gibs_11_reset = reset;
  assign gibs_11_io_cfg_en = cfgRegs_3[44]; // @[CGRA.scala 509:38]
  assign gibs_11_io_cfg_addr = cfgRegs_3[43:32]; // @[CGRA.scala 510:38]
  assign gibs_11_io_cfg_data = cfgRegs_3[31:0]; // @[CGRA.scala 511:38]
  assign gibs_11_io_opinNW_0 = pes_1_io_out_0; // @[CGRA.scala 401:47]
  assign gibs_11_io_opinNE_0 = pes_2_io_out_0; // @[CGRA.scala 400:45]
  assign gibs_11_io_opinSE_0 = pes_10_io_out_0; // @[CGRA.scala 398:41]
  assign gibs_11_io_opinSW_0 = pes_9_io_out_0; // @[CGRA.scala 399:43]
  assign gibs_11_io_itrackW_0 = gibs_10_io_otrackE_0; // @[CGRA.scala 466:16]
  assign gibs_11_io_itrackN_0 = gibs_2_io_otrackS_0; // @[CGRA.scala 436:16]
  assign gibs_11_io_itrackE_0 = gibs_12_io_otrackW_0; // @[CGRA.scala 472:16]
  assign gibs_11_io_itrackS_0 = gibs_20_io_otrackN_0; // @[CGRA.scala 442:16]
  assign gibs_12_clock = clock;
  assign gibs_12_reset = reset;
  assign gibs_12_io_cfg_en = cfgRegs_3[44]; // @[CGRA.scala 509:38]
  assign gibs_12_io_cfg_addr = cfgRegs_3[43:32]; // @[CGRA.scala 510:38]
  assign gibs_12_io_cfg_data = cfgRegs_3[31:0]; // @[CGRA.scala 511:38]
  assign gibs_12_io_opinNW_0 = pes_2_io_out_0; // @[CGRA.scala 401:47]
  assign gibs_12_io_opinNE_0 = pes_3_io_out_0; // @[CGRA.scala 400:45]
  assign gibs_12_io_opinSE_0 = pes_11_io_out_0; // @[CGRA.scala 398:41]
  assign gibs_12_io_opinSW_0 = pes_10_io_out_0; // @[CGRA.scala 399:43]
  assign gibs_12_io_itrackW_0 = gibs_11_io_otrackE_0; // @[CGRA.scala 466:16]
  assign gibs_12_io_itrackN_0 = gibs_3_io_otrackS_0; // @[CGRA.scala 436:16]
  assign gibs_12_io_itrackE_0 = gibs_13_io_otrackW_0; // @[CGRA.scala 472:16]
  assign gibs_12_io_itrackS_0 = gibs_21_io_otrackN_0; // @[CGRA.scala 442:16]
  assign gibs_13_clock = clock;
  assign gibs_13_reset = reset;
  assign gibs_13_io_cfg_en = cfgRegs_3[44]; // @[CGRA.scala 509:38]
  assign gibs_13_io_cfg_addr = cfgRegs_3[43:32]; // @[CGRA.scala 510:38]
  assign gibs_13_io_cfg_data = cfgRegs_3[31:0]; // @[CGRA.scala 511:38]
  assign gibs_13_io_opinNW_0 = pes_3_io_out_0; // @[CGRA.scala 401:47]
  assign gibs_13_io_opinNE_0 = pes_4_io_out_0; // @[CGRA.scala 400:45]
  assign gibs_13_io_opinSE_0 = pes_12_io_out_0; // @[CGRA.scala 398:41]
  assign gibs_13_io_opinSW_0 = pes_11_io_out_0; // @[CGRA.scala 399:43]
  assign gibs_13_io_itrackW_0 = gibs_12_io_otrackE_0; // @[CGRA.scala 466:16]
  assign gibs_13_io_itrackN_0 = gibs_4_io_otrackS_0; // @[CGRA.scala 436:16]
  assign gibs_13_io_itrackE_0 = gibs_14_io_otrackW_0; // @[CGRA.scala 472:16]
  assign gibs_13_io_itrackS_0 = gibs_22_io_otrackN_0; // @[CGRA.scala 442:16]
  assign gibs_14_clock = clock;
  assign gibs_14_reset = reset;
  assign gibs_14_io_cfg_en = cfgRegs_3[44]; // @[CGRA.scala 509:38]
  assign gibs_14_io_cfg_addr = cfgRegs_3[43:32]; // @[CGRA.scala 510:38]
  assign gibs_14_io_cfg_data = cfgRegs_3[31:0]; // @[CGRA.scala 511:38]
  assign gibs_14_io_opinNW_0 = pes_4_io_out_0; // @[CGRA.scala 401:47]
  assign gibs_14_io_opinNE_0 = pes_5_io_out_0; // @[CGRA.scala 400:45]
  assign gibs_14_io_opinSE_0 = pes_13_io_out_0; // @[CGRA.scala 398:41]
  assign gibs_14_io_opinSW_0 = pes_12_io_out_0; // @[CGRA.scala 399:43]
  assign gibs_14_io_itrackW_0 = gibs_13_io_otrackE_0; // @[CGRA.scala 466:16]
  assign gibs_14_io_itrackN_0 = gibs_5_io_otrackS_0; // @[CGRA.scala 436:16]
  assign gibs_14_io_itrackE_0 = gibs_15_io_otrackW_0; // @[CGRA.scala 472:16]
  assign gibs_14_io_itrackS_0 = gibs_23_io_otrackN_0; // @[CGRA.scala 442:16]
  assign gibs_15_clock = clock;
  assign gibs_15_reset = reset;
  assign gibs_15_io_cfg_en = cfgRegs_3[44]; // @[CGRA.scala 509:38]
  assign gibs_15_io_cfg_addr = cfgRegs_3[43:32]; // @[CGRA.scala 510:38]
  assign gibs_15_io_cfg_data = cfgRegs_3[31:0]; // @[CGRA.scala 511:38]
  assign gibs_15_io_opinNW_0 = pes_5_io_out_0; // @[CGRA.scala 401:47]
  assign gibs_15_io_opinNE_0 = pes_6_io_out_0; // @[CGRA.scala 400:45]
  assign gibs_15_io_opinSE_0 = pes_14_io_out_0; // @[CGRA.scala 398:41]
  assign gibs_15_io_opinSW_0 = pes_13_io_out_0; // @[CGRA.scala 399:43]
  assign gibs_15_io_itrackW_0 = gibs_14_io_otrackE_0; // @[CGRA.scala 466:16]
  assign gibs_15_io_itrackN_0 = gibs_6_io_otrackS_0; // @[CGRA.scala 436:16]
  assign gibs_15_io_itrackE_0 = gibs_16_io_otrackW_0; // @[CGRA.scala 472:16]
  assign gibs_15_io_itrackS_0 = gibs_24_io_otrackN_0; // @[CGRA.scala 442:16]
  assign gibs_16_clock = clock;
  assign gibs_16_reset = reset;
  assign gibs_16_io_cfg_en = cfgRegs_3[44]; // @[CGRA.scala 509:38]
  assign gibs_16_io_cfg_addr = cfgRegs_3[43:32]; // @[CGRA.scala 510:38]
  assign gibs_16_io_cfg_data = cfgRegs_3[31:0]; // @[CGRA.scala 511:38]
  assign gibs_16_io_opinNW_0 = pes_6_io_out_0; // @[CGRA.scala 401:47]
  assign gibs_16_io_opinNE_0 = pes_7_io_out_0; // @[CGRA.scala 400:45]
  assign gibs_16_io_opinSE_0 = pes_15_io_out_0; // @[CGRA.scala 398:41]
  assign gibs_16_io_opinSW_0 = pes_14_io_out_0; // @[CGRA.scala 399:43]
  assign gibs_16_io_itrackW_0 = gibs_15_io_otrackE_0; // @[CGRA.scala 466:16]
  assign gibs_16_io_itrackN_0 = gibs_7_io_otrackS_0; // @[CGRA.scala 436:16]
  assign gibs_16_io_itrackE_0 = gibs_17_io_otrackW_0; // @[CGRA.scala 472:16]
  assign gibs_16_io_itrackS_0 = gibs_25_io_otrackN_0; // @[CGRA.scala 442:16]
  assign gibs_17_clock = clock;
  assign gibs_17_reset = reset;
  assign gibs_17_io_cfg_en = cfgRegs_3[44]; // @[CGRA.scala 509:38]
  assign gibs_17_io_cfg_addr = cfgRegs_3[43:32]; // @[CGRA.scala 510:38]
  assign gibs_17_io_cfg_data = cfgRegs_3[31:0]; // @[CGRA.scala 511:38]
  assign gibs_17_io_opinNW_0 = pes_7_io_out_0; // @[CGRA.scala 401:47]
  assign gibs_17_io_opinSW_0 = pes_15_io_out_0; // @[CGRA.scala 399:43]
  assign gibs_17_io_itrackW_0 = gibs_16_io_otrackE_0; // @[CGRA.scala 459:16]
  assign gibs_17_io_itrackN_0 = gibs_8_io_otrackS_0; // @[CGRA.scala 436:16]
  assign gibs_17_io_itrackS_0 = gibs_26_io_otrackN_0; // @[CGRA.scala 442:16]
  assign gibs_18_clock = clock;
  assign gibs_18_reset = reset;
  assign gibs_18_io_cfg_en = cfgRegs_5[44]; // @[CGRA.scala 509:38]
  assign gibs_18_io_cfg_addr = cfgRegs_5[43:32]; // @[CGRA.scala 510:38]
  assign gibs_18_io_cfg_data = cfgRegs_5[31:0]; // @[CGRA.scala 511:38]
  assign gibs_18_io_opinNE_0 = pes_8_io_out_0; // @[CGRA.scala 400:45]
  assign gibs_18_io_opinSE_0 = pes_16_io_out_0; // @[CGRA.scala 398:41]
  assign gibs_18_io_itrackN_0 = gibs_9_io_otrackS_0; // @[CGRA.scala 436:16]
  assign gibs_18_io_itrackE_0 = gibs_19_io_otrackW_0; // @[CGRA.scala 451:16]
  assign gibs_18_io_itrackS_0 = gibs_27_io_otrackN_0; // @[CGRA.scala 442:16]
  assign gibs_19_clock = clock;
  assign gibs_19_reset = reset;
  assign gibs_19_io_cfg_en = cfgRegs_5[44]; // @[CGRA.scala 509:38]
  assign gibs_19_io_cfg_addr = cfgRegs_5[43:32]; // @[CGRA.scala 510:38]
  assign gibs_19_io_cfg_data = cfgRegs_5[31:0]; // @[CGRA.scala 511:38]
  assign gibs_19_io_opinNW_0 = pes_8_io_out_0; // @[CGRA.scala 401:47]
  assign gibs_19_io_opinNE_0 = pes_9_io_out_0; // @[CGRA.scala 400:45]
  assign gibs_19_io_opinSE_0 = pes_17_io_out_0; // @[CGRA.scala 398:41]
  assign gibs_19_io_opinSW_0 = pes_16_io_out_0; // @[CGRA.scala 399:43]
  assign gibs_19_io_itrackW_0 = gibs_18_io_otrackE_0; // @[CGRA.scala 466:16]
  assign gibs_19_io_itrackN_0 = gibs_10_io_otrackS_0; // @[CGRA.scala 436:16]
  assign gibs_19_io_itrackE_0 = gibs_20_io_otrackW_0; // @[CGRA.scala 472:16]
  assign gibs_19_io_itrackS_0 = gibs_28_io_otrackN_0; // @[CGRA.scala 442:16]
  assign gibs_20_clock = clock;
  assign gibs_20_reset = reset;
  assign gibs_20_io_cfg_en = cfgRegs_5[44]; // @[CGRA.scala 509:38]
  assign gibs_20_io_cfg_addr = cfgRegs_5[43:32]; // @[CGRA.scala 510:38]
  assign gibs_20_io_cfg_data = cfgRegs_5[31:0]; // @[CGRA.scala 511:38]
  assign gibs_20_io_opinNW_0 = pes_9_io_out_0; // @[CGRA.scala 401:47]
  assign gibs_20_io_opinNE_0 = pes_10_io_out_0; // @[CGRA.scala 400:45]
  assign gibs_20_io_opinSE_0 = pes_18_io_out_0; // @[CGRA.scala 398:41]
  assign gibs_20_io_opinSW_0 = pes_17_io_out_0; // @[CGRA.scala 399:43]
  assign gibs_20_io_itrackW_0 = gibs_19_io_otrackE_0; // @[CGRA.scala 466:16]
  assign gibs_20_io_itrackN_0 = gibs_11_io_otrackS_0; // @[CGRA.scala 436:16]
  assign gibs_20_io_itrackE_0 = gibs_21_io_otrackW_0; // @[CGRA.scala 472:16]
  assign gibs_20_io_itrackS_0 = gibs_29_io_otrackN_0; // @[CGRA.scala 442:16]
  assign gibs_21_clock = clock;
  assign gibs_21_reset = reset;
  assign gibs_21_io_cfg_en = cfgRegs_5[44]; // @[CGRA.scala 509:38]
  assign gibs_21_io_cfg_addr = cfgRegs_5[43:32]; // @[CGRA.scala 510:38]
  assign gibs_21_io_cfg_data = cfgRegs_5[31:0]; // @[CGRA.scala 511:38]
  assign gibs_21_io_opinNW_0 = pes_10_io_out_0; // @[CGRA.scala 401:47]
  assign gibs_21_io_opinNE_0 = pes_11_io_out_0; // @[CGRA.scala 400:45]
  assign gibs_21_io_opinSE_0 = pes_19_io_out_0; // @[CGRA.scala 398:41]
  assign gibs_21_io_opinSW_0 = pes_18_io_out_0; // @[CGRA.scala 399:43]
  assign gibs_21_io_itrackW_0 = gibs_20_io_otrackE_0; // @[CGRA.scala 466:16]
  assign gibs_21_io_itrackN_0 = gibs_12_io_otrackS_0; // @[CGRA.scala 436:16]
  assign gibs_21_io_itrackE_0 = gibs_22_io_otrackW_0; // @[CGRA.scala 472:16]
  assign gibs_21_io_itrackS_0 = gibs_30_io_otrackN_0; // @[CGRA.scala 442:16]
  assign gibs_22_clock = clock;
  assign gibs_22_reset = reset;
  assign gibs_22_io_cfg_en = cfgRegs_5[44]; // @[CGRA.scala 509:38]
  assign gibs_22_io_cfg_addr = cfgRegs_5[43:32]; // @[CGRA.scala 510:38]
  assign gibs_22_io_cfg_data = cfgRegs_5[31:0]; // @[CGRA.scala 511:38]
  assign gibs_22_io_opinNW_0 = pes_11_io_out_0; // @[CGRA.scala 401:47]
  assign gibs_22_io_opinNE_0 = pes_12_io_out_0; // @[CGRA.scala 400:45]
  assign gibs_22_io_opinSE_0 = pes_20_io_out_0; // @[CGRA.scala 398:41]
  assign gibs_22_io_opinSW_0 = pes_19_io_out_0; // @[CGRA.scala 399:43]
  assign gibs_22_io_itrackW_0 = gibs_21_io_otrackE_0; // @[CGRA.scala 466:16]
  assign gibs_22_io_itrackN_0 = gibs_13_io_otrackS_0; // @[CGRA.scala 436:16]
  assign gibs_22_io_itrackE_0 = gibs_23_io_otrackW_0; // @[CGRA.scala 472:16]
  assign gibs_22_io_itrackS_0 = gibs_31_io_otrackN_0; // @[CGRA.scala 442:16]
  assign gibs_23_clock = clock;
  assign gibs_23_reset = reset;
  assign gibs_23_io_cfg_en = cfgRegs_5[44]; // @[CGRA.scala 509:38]
  assign gibs_23_io_cfg_addr = cfgRegs_5[43:32]; // @[CGRA.scala 510:38]
  assign gibs_23_io_cfg_data = cfgRegs_5[31:0]; // @[CGRA.scala 511:38]
  assign gibs_23_io_opinNW_0 = pes_12_io_out_0; // @[CGRA.scala 401:47]
  assign gibs_23_io_opinNE_0 = pes_13_io_out_0; // @[CGRA.scala 400:45]
  assign gibs_23_io_opinSE_0 = pes_21_io_out_0; // @[CGRA.scala 398:41]
  assign gibs_23_io_opinSW_0 = pes_20_io_out_0; // @[CGRA.scala 399:43]
  assign gibs_23_io_itrackW_0 = gibs_22_io_otrackE_0; // @[CGRA.scala 466:16]
  assign gibs_23_io_itrackN_0 = gibs_14_io_otrackS_0; // @[CGRA.scala 436:16]
  assign gibs_23_io_itrackE_0 = gibs_24_io_otrackW_0; // @[CGRA.scala 472:16]
  assign gibs_23_io_itrackS_0 = gibs_32_io_otrackN_0; // @[CGRA.scala 442:16]
  assign gibs_24_clock = clock;
  assign gibs_24_reset = reset;
  assign gibs_24_io_cfg_en = cfgRegs_5[44]; // @[CGRA.scala 509:38]
  assign gibs_24_io_cfg_addr = cfgRegs_5[43:32]; // @[CGRA.scala 510:38]
  assign gibs_24_io_cfg_data = cfgRegs_5[31:0]; // @[CGRA.scala 511:38]
  assign gibs_24_io_opinNW_0 = pes_13_io_out_0; // @[CGRA.scala 401:47]
  assign gibs_24_io_opinNE_0 = pes_14_io_out_0; // @[CGRA.scala 400:45]
  assign gibs_24_io_opinSE_0 = pes_22_io_out_0; // @[CGRA.scala 398:41]
  assign gibs_24_io_opinSW_0 = pes_21_io_out_0; // @[CGRA.scala 399:43]
  assign gibs_24_io_itrackW_0 = gibs_23_io_otrackE_0; // @[CGRA.scala 466:16]
  assign gibs_24_io_itrackN_0 = gibs_15_io_otrackS_0; // @[CGRA.scala 436:16]
  assign gibs_24_io_itrackE_0 = gibs_25_io_otrackW_0; // @[CGRA.scala 472:16]
  assign gibs_24_io_itrackS_0 = gibs_33_io_otrackN_0; // @[CGRA.scala 442:16]
  assign gibs_25_clock = clock;
  assign gibs_25_reset = reset;
  assign gibs_25_io_cfg_en = cfgRegs_5[44]; // @[CGRA.scala 509:38]
  assign gibs_25_io_cfg_addr = cfgRegs_5[43:32]; // @[CGRA.scala 510:38]
  assign gibs_25_io_cfg_data = cfgRegs_5[31:0]; // @[CGRA.scala 511:38]
  assign gibs_25_io_opinNW_0 = pes_14_io_out_0; // @[CGRA.scala 401:47]
  assign gibs_25_io_opinNE_0 = pes_15_io_out_0; // @[CGRA.scala 400:45]
  assign gibs_25_io_opinSE_0 = pes_23_io_out_0; // @[CGRA.scala 398:41]
  assign gibs_25_io_opinSW_0 = pes_22_io_out_0; // @[CGRA.scala 399:43]
  assign gibs_25_io_itrackW_0 = gibs_24_io_otrackE_0; // @[CGRA.scala 466:16]
  assign gibs_25_io_itrackN_0 = gibs_16_io_otrackS_0; // @[CGRA.scala 436:16]
  assign gibs_25_io_itrackE_0 = gibs_26_io_otrackW_0; // @[CGRA.scala 472:16]
  assign gibs_25_io_itrackS_0 = gibs_34_io_otrackN_0; // @[CGRA.scala 442:16]
  assign gibs_26_clock = clock;
  assign gibs_26_reset = reset;
  assign gibs_26_io_cfg_en = cfgRegs_5[44]; // @[CGRA.scala 509:38]
  assign gibs_26_io_cfg_addr = cfgRegs_5[43:32]; // @[CGRA.scala 510:38]
  assign gibs_26_io_cfg_data = cfgRegs_5[31:0]; // @[CGRA.scala 511:38]
  assign gibs_26_io_opinNW_0 = pes_15_io_out_0; // @[CGRA.scala 401:47]
  assign gibs_26_io_opinSW_0 = pes_23_io_out_0; // @[CGRA.scala 399:43]
  assign gibs_26_io_itrackW_0 = gibs_25_io_otrackE_0; // @[CGRA.scala 459:16]
  assign gibs_26_io_itrackN_0 = gibs_17_io_otrackS_0; // @[CGRA.scala 436:16]
  assign gibs_26_io_itrackS_0 = gibs_35_io_otrackN_0; // @[CGRA.scala 442:16]
  assign gibs_27_clock = clock;
  assign gibs_27_reset = reset;
  assign gibs_27_io_cfg_en = cfgRegs_7[44]; // @[CGRA.scala 509:38]
  assign gibs_27_io_cfg_addr = cfgRegs_7[43:32]; // @[CGRA.scala 510:38]
  assign gibs_27_io_cfg_data = cfgRegs_7[31:0]; // @[CGRA.scala 511:38]
  assign gibs_27_io_opinNE_0 = pes_16_io_out_0; // @[CGRA.scala 400:45]
  assign gibs_27_io_opinSE_0 = pes_24_io_out_0; // @[CGRA.scala 398:41]
  assign gibs_27_io_itrackN_0 = gibs_18_io_otrackS_0; // @[CGRA.scala 436:16]
  assign gibs_27_io_itrackE_0 = gibs_28_io_otrackW_0; // @[CGRA.scala 451:16]
  assign gibs_27_io_itrackS_0 = gibs_36_io_otrackN_0; // @[CGRA.scala 442:16]
  assign gibs_28_clock = clock;
  assign gibs_28_reset = reset;
  assign gibs_28_io_cfg_en = cfgRegs_7[44]; // @[CGRA.scala 509:38]
  assign gibs_28_io_cfg_addr = cfgRegs_7[43:32]; // @[CGRA.scala 510:38]
  assign gibs_28_io_cfg_data = cfgRegs_7[31:0]; // @[CGRA.scala 511:38]
  assign gibs_28_io_opinNW_0 = pes_16_io_out_0; // @[CGRA.scala 401:47]
  assign gibs_28_io_opinNE_0 = pes_17_io_out_0; // @[CGRA.scala 400:45]
  assign gibs_28_io_opinSE_0 = pes_25_io_out_0; // @[CGRA.scala 398:41]
  assign gibs_28_io_opinSW_0 = pes_24_io_out_0; // @[CGRA.scala 399:43]
  assign gibs_28_io_itrackW_0 = gibs_27_io_otrackE_0; // @[CGRA.scala 466:16]
  assign gibs_28_io_itrackN_0 = gibs_19_io_otrackS_0; // @[CGRA.scala 436:16]
  assign gibs_28_io_itrackE_0 = gibs_29_io_otrackW_0; // @[CGRA.scala 472:16]
  assign gibs_28_io_itrackS_0 = gibs_37_io_otrackN_0; // @[CGRA.scala 442:16]
  assign gibs_29_clock = clock;
  assign gibs_29_reset = reset;
  assign gibs_29_io_cfg_en = cfgRegs_7[44]; // @[CGRA.scala 509:38]
  assign gibs_29_io_cfg_addr = cfgRegs_7[43:32]; // @[CGRA.scala 510:38]
  assign gibs_29_io_cfg_data = cfgRegs_7[31:0]; // @[CGRA.scala 511:38]
  assign gibs_29_io_opinNW_0 = pes_17_io_out_0; // @[CGRA.scala 401:47]
  assign gibs_29_io_opinNE_0 = pes_18_io_out_0; // @[CGRA.scala 400:45]
  assign gibs_29_io_opinSE_0 = pes_26_io_out_0; // @[CGRA.scala 398:41]
  assign gibs_29_io_opinSW_0 = pes_25_io_out_0; // @[CGRA.scala 399:43]
  assign gibs_29_io_itrackW_0 = gibs_28_io_otrackE_0; // @[CGRA.scala 466:16]
  assign gibs_29_io_itrackN_0 = gibs_20_io_otrackS_0; // @[CGRA.scala 436:16]
  assign gibs_29_io_itrackE_0 = gibs_30_io_otrackW_0; // @[CGRA.scala 472:16]
  assign gibs_29_io_itrackS_0 = gibs_38_io_otrackN_0; // @[CGRA.scala 442:16]
  assign gibs_30_clock = clock;
  assign gibs_30_reset = reset;
  assign gibs_30_io_cfg_en = cfgRegs_7[44]; // @[CGRA.scala 509:38]
  assign gibs_30_io_cfg_addr = cfgRegs_7[43:32]; // @[CGRA.scala 510:38]
  assign gibs_30_io_cfg_data = cfgRegs_7[31:0]; // @[CGRA.scala 511:38]
  assign gibs_30_io_opinNW_0 = pes_18_io_out_0; // @[CGRA.scala 401:47]
  assign gibs_30_io_opinNE_0 = pes_19_io_out_0; // @[CGRA.scala 400:45]
  assign gibs_30_io_opinSE_0 = pes_27_io_out_0; // @[CGRA.scala 398:41]
  assign gibs_30_io_opinSW_0 = pes_26_io_out_0; // @[CGRA.scala 399:43]
  assign gibs_30_io_itrackW_0 = gibs_29_io_otrackE_0; // @[CGRA.scala 466:16]
  assign gibs_30_io_itrackN_0 = gibs_21_io_otrackS_0; // @[CGRA.scala 436:16]
  assign gibs_30_io_itrackE_0 = gibs_31_io_otrackW_0; // @[CGRA.scala 472:16]
  assign gibs_30_io_itrackS_0 = gibs_39_io_otrackN_0; // @[CGRA.scala 442:16]
  assign gibs_31_clock = clock;
  assign gibs_31_reset = reset;
  assign gibs_31_io_cfg_en = cfgRegs_7[44]; // @[CGRA.scala 509:38]
  assign gibs_31_io_cfg_addr = cfgRegs_7[43:32]; // @[CGRA.scala 510:38]
  assign gibs_31_io_cfg_data = cfgRegs_7[31:0]; // @[CGRA.scala 511:38]
  assign gibs_31_io_opinNW_0 = pes_19_io_out_0; // @[CGRA.scala 401:47]
  assign gibs_31_io_opinNE_0 = pes_20_io_out_0; // @[CGRA.scala 400:45]
  assign gibs_31_io_opinSE_0 = pes_28_io_out_0; // @[CGRA.scala 398:41]
  assign gibs_31_io_opinSW_0 = pes_27_io_out_0; // @[CGRA.scala 399:43]
  assign gibs_31_io_itrackW_0 = gibs_30_io_otrackE_0; // @[CGRA.scala 466:16]
  assign gibs_31_io_itrackN_0 = gibs_22_io_otrackS_0; // @[CGRA.scala 436:16]
  assign gibs_31_io_itrackE_0 = gibs_32_io_otrackW_0; // @[CGRA.scala 472:16]
  assign gibs_31_io_itrackS_0 = gibs_40_io_otrackN_0; // @[CGRA.scala 442:16]
  assign gibs_32_clock = clock;
  assign gibs_32_reset = reset;
  assign gibs_32_io_cfg_en = cfgRegs_7[44]; // @[CGRA.scala 509:38]
  assign gibs_32_io_cfg_addr = cfgRegs_7[43:32]; // @[CGRA.scala 510:38]
  assign gibs_32_io_cfg_data = cfgRegs_7[31:0]; // @[CGRA.scala 511:38]
  assign gibs_32_io_opinNW_0 = pes_20_io_out_0; // @[CGRA.scala 401:47]
  assign gibs_32_io_opinNE_0 = pes_21_io_out_0; // @[CGRA.scala 400:45]
  assign gibs_32_io_opinSE_0 = pes_29_io_out_0; // @[CGRA.scala 398:41]
  assign gibs_32_io_opinSW_0 = pes_28_io_out_0; // @[CGRA.scala 399:43]
  assign gibs_32_io_itrackW_0 = gibs_31_io_otrackE_0; // @[CGRA.scala 466:16]
  assign gibs_32_io_itrackN_0 = gibs_23_io_otrackS_0; // @[CGRA.scala 436:16]
  assign gibs_32_io_itrackE_0 = gibs_33_io_otrackW_0; // @[CGRA.scala 472:16]
  assign gibs_32_io_itrackS_0 = gibs_41_io_otrackN_0; // @[CGRA.scala 442:16]
  assign gibs_33_clock = clock;
  assign gibs_33_reset = reset;
  assign gibs_33_io_cfg_en = cfgRegs_7[44]; // @[CGRA.scala 509:38]
  assign gibs_33_io_cfg_addr = cfgRegs_7[43:32]; // @[CGRA.scala 510:38]
  assign gibs_33_io_cfg_data = cfgRegs_7[31:0]; // @[CGRA.scala 511:38]
  assign gibs_33_io_opinNW_0 = pes_21_io_out_0; // @[CGRA.scala 401:47]
  assign gibs_33_io_opinNE_0 = pes_22_io_out_0; // @[CGRA.scala 400:45]
  assign gibs_33_io_opinSE_0 = pes_30_io_out_0; // @[CGRA.scala 398:41]
  assign gibs_33_io_opinSW_0 = pes_29_io_out_0; // @[CGRA.scala 399:43]
  assign gibs_33_io_itrackW_0 = gibs_32_io_otrackE_0; // @[CGRA.scala 466:16]
  assign gibs_33_io_itrackN_0 = gibs_24_io_otrackS_0; // @[CGRA.scala 436:16]
  assign gibs_33_io_itrackE_0 = gibs_34_io_otrackW_0; // @[CGRA.scala 472:16]
  assign gibs_33_io_itrackS_0 = gibs_42_io_otrackN_0; // @[CGRA.scala 442:16]
  assign gibs_34_clock = clock;
  assign gibs_34_reset = reset;
  assign gibs_34_io_cfg_en = cfgRegs_7[44]; // @[CGRA.scala 509:38]
  assign gibs_34_io_cfg_addr = cfgRegs_7[43:32]; // @[CGRA.scala 510:38]
  assign gibs_34_io_cfg_data = cfgRegs_7[31:0]; // @[CGRA.scala 511:38]
  assign gibs_34_io_opinNW_0 = pes_22_io_out_0; // @[CGRA.scala 401:47]
  assign gibs_34_io_opinNE_0 = pes_23_io_out_0; // @[CGRA.scala 400:45]
  assign gibs_34_io_opinSE_0 = pes_31_io_out_0; // @[CGRA.scala 398:41]
  assign gibs_34_io_opinSW_0 = pes_30_io_out_0; // @[CGRA.scala 399:43]
  assign gibs_34_io_itrackW_0 = gibs_33_io_otrackE_0; // @[CGRA.scala 466:16]
  assign gibs_34_io_itrackN_0 = gibs_25_io_otrackS_0; // @[CGRA.scala 436:16]
  assign gibs_34_io_itrackE_0 = gibs_35_io_otrackW_0; // @[CGRA.scala 472:16]
  assign gibs_34_io_itrackS_0 = gibs_43_io_otrackN_0; // @[CGRA.scala 442:16]
  assign gibs_35_clock = clock;
  assign gibs_35_reset = reset;
  assign gibs_35_io_cfg_en = cfgRegs_7[44]; // @[CGRA.scala 509:38]
  assign gibs_35_io_cfg_addr = cfgRegs_7[43:32]; // @[CGRA.scala 510:38]
  assign gibs_35_io_cfg_data = cfgRegs_7[31:0]; // @[CGRA.scala 511:38]
  assign gibs_35_io_opinNW_0 = pes_23_io_out_0; // @[CGRA.scala 401:47]
  assign gibs_35_io_opinSW_0 = pes_31_io_out_0; // @[CGRA.scala 399:43]
  assign gibs_35_io_itrackW_0 = gibs_34_io_otrackE_0; // @[CGRA.scala 459:16]
  assign gibs_35_io_itrackN_0 = gibs_26_io_otrackS_0; // @[CGRA.scala 436:16]
  assign gibs_35_io_itrackS_0 = gibs_44_io_otrackN_0; // @[CGRA.scala 442:16]
  assign gibs_36_clock = clock;
  assign gibs_36_reset = reset;
  assign gibs_36_io_cfg_en = cfgRegs_9[44]; // @[CGRA.scala 509:38]
  assign gibs_36_io_cfg_addr = cfgRegs_9[43:32]; // @[CGRA.scala 510:38]
  assign gibs_36_io_cfg_data = cfgRegs_9[31:0]; // @[CGRA.scala 511:38]
  assign gibs_36_io_opinNE_0 = pes_24_io_out_0; // @[CGRA.scala 400:45]
  assign gibs_36_io_opinSE_0 = pes_32_io_out_0; // @[CGRA.scala 398:41]
  assign gibs_36_io_itrackN_0 = gibs_27_io_otrackS_0; // @[CGRA.scala 436:16]
  assign gibs_36_io_itrackE_0 = gibs_37_io_otrackW_0; // @[CGRA.scala 451:16]
  assign gibs_36_io_itrackS_0 = gibs_45_io_otrackN_0; // @[CGRA.scala 442:16]
  assign gibs_37_clock = clock;
  assign gibs_37_reset = reset;
  assign gibs_37_io_cfg_en = cfgRegs_9[44]; // @[CGRA.scala 509:38]
  assign gibs_37_io_cfg_addr = cfgRegs_9[43:32]; // @[CGRA.scala 510:38]
  assign gibs_37_io_cfg_data = cfgRegs_9[31:0]; // @[CGRA.scala 511:38]
  assign gibs_37_io_opinNW_0 = pes_24_io_out_0; // @[CGRA.scala 401:47]
  assign gibs_37_io_opinNE_0 = pes_25_io_out_0; // @[CGRA.scala 400:45]
  assign gibs_37_io_opinSE_0 = pes_33_io_out_0; // @[CGRA.scala 398:41]
  assign gibs_37_io_opinSW_0 = pes_32_io_out_0; // @[CGRA.scala 399:43]
  assign gibs_37_io_itrackW_0 = gibs_36_io_otrackE_0; // @[CGRA.scala 466:16]
  assign gibs_37_io_itrackN_0 = gibs_28_io_otrackS_0; // @[CGRA.scala 436:16]
  assign gibs_37_io_itrackE_0 = gibs_38_io_otrackW_0; // @[CGRA.scala 472:16]
  assign gibs_37_io_itrackS_0 = gibs_46_io_otrackN_0; // @[CGRA.scala 442:16]
  assign gibs_38_clock = clock;
  assign gibs_38_reset = reset;
  assign gibs_38_io_cfg_en = cfgRegs_9[44]; // @[CGRA.scala 509:38]
  assign gibs_38_io_cfg_addr = cfgRegs_9[43:32]; // @[CGRA.scala 510:38]
  assign gibs_38_io_cfg_data = cfgRegs_9[31:0]; // @[CGRA.scala 511:38]
  assign gibs_38_io_opinNW_0 = pes_25_io_out_0; // @[CGRA.scala 401:47]
  assign gibs_38_io_opinNE_0 = pes_26_io_out_0; // @[CGRA.scala 400:45]
  assign gibs_38_io_opinSE_0 = pes_34_io_out_0; // @[CGRA.scala 398:41]
  assign gibs_38_io_opinSW_0 = pes_33_io_out_0; // @[CGRA.scala 399:43]
  assign gibs_38_io_itrackW_0 = gibs_37_io_otrackE_0; // @[CGRA.scala 466:16]
  assign gibs_38_io_itrackN_0 = gibs_29_io_otrackS_0; // @[CGRA.scala 436:16]
  assign gibs_38_io_itrackE_0 = gibs_39_io_otrackW_0; // @[CGRA.scala 472:16]
  assign gibs_38_io_itrackS_0 = gibs_47_io_otrackN_0; // @[CGRA.scala 442:16]
  assign gibs_39_clock = clock;
  assign gibs_39_reset = reset;
  assign gibs_39_io_cfg_en = cfgRegs_9[44]; // @[CGRA.scala 509:38]
  assign gibs_39_io_cfg_addr = cfgRegs_9[43:32]; // @[CGRA.scala 510:38]
  assign gibs_39_io_cfg_data = cfgRegs_9[31:0]; // @[CGRA.scala 511:38]
  assign gibs_39_io_opinNW_0 = pes_26_io_out_0; // @[CGRA.scala 401:47]
  assign gibs_39_io_opinNE_0 = pes_27_io_out_0; // @[CGRA.scala 400:45]
  assign gibs_39_io_opinSE_0 = pes_35_io_out_0; // @[CGRA.scala 398:41]
  assign gibs_39_io_opinSW_0 = pes_34_io_out_0; // @[CGRA.scala 399:43]
  assign gibs_39_io_itrackW_0 = gibs_38_io_otrackE_0; // @[CGRA.scala 466:16]
  assign gibs_39_io_itrackN_0 = gibs_30_io_otrackS_0; // @[CGRA.scala 436:16]
  assign gibs_39_io_itrackE_0 = gibs_40_io_otrackW_0; // @[CGRA.scala 472:16]
  assign gibs_39_io_itrackS_0 = gibs_48_io_otrackN_0; // @[CGRA.scala 442:16]
  assign gibs_40_clock = clock;
  assign gibs_40_reset = reset;
  assign gibs_40_io_cfg_en = cfgRegs_9[44]; // @[CGRA.scala 509:38]
  assign gibs_40_io_cfg_addr = cfgRegs_9[43:32]; // @[CGRA.scala 510:38]
  assign gibs_40_io_cfg_data = cfgRegs_9[31:0]; // @[CGRA.scala 511:38]
  assign gibs_40_io_opinNW_0 = pes_27_io_out_0; // @[CGRA.scala 401:47]
  assign gibs_40_io_opinNE_0 = pes_28_io_out_0; // @[CGRA.scala 400:45]
  assign gibs_40_io_opinSE_0 = pes_36_io_out_0; // @[CGRA.scala 398:41]
  assign gibs_40_io_opinSW_0 = pes_35_io_out_0; // @[CGRA.scala 399:43]
  assign gibs_40_io_itrackW_0 = gibs_39_io_otrackE_0; // @[CGRA.scala 466:16]
  assign gibs_40_io_itrackN_0 = gibs_31_io_otrackS_0; // @[CGRA.scala 436:16]
  assign gibs_40_io_itrackE_0 = gibs_41_io_otrackW_0; // @[CGRA.scala 472:16]
  assign gibs_40_io_itrackS_0 = gibs_49_io_otrackN_0; // @[CGRA.scala 442:16]
  assign gibs_41_clock = clock;
  assign gibs_41_reset = reset;
  assign gibs_41_io_cfg_en = cfgRegs_9[44]; // @[CGRA.scala 509:38]
  assign gibs_41_io_cfg_addr = cfgRegs_9[43:32]; // @[CGRA.scala 510:38]
  assign gibs_41_io_cfg_data = cfgRegs_9[31:0]; // @[CGRA.scala 511:38]
  assign gibs_41_io_opinNW_0 = pes_28_io_out_0; // @[CGRA.scala 401:47]
  assign gibs_41_io_opinNE_0 = pes_29_io_out_0; // @[CGRA.scala 400:45]
  assign gibs_41_io_opinSE_0 = pes_37_io_out_0; // @[CGRA.scala 398:41]
  assign gibs_41_io_opinSW_0 = pes_36_io_out_0; // @[CGRA.scala 399:43]
  assign gibs_41_io_itrackW_0 = gibs_40_io_otrackE_0; // @[CGRA.scala 466:16]
  assign gibs_41_io_itrackN_0 = gibs_32_io_otrackS_0; // @[CGRA.scala 436:16]
  assign gibs_41_io_itrackE_0 = gibs_42_io_otrackW_0; // @[CGRA.scala 472:16]
  assign gibs_41_io_itrackS_0 = gibs_50_io_otrackN_0; // @[CGRA.scala 442:16]
  assign gibs_42_clock = clock;
  assign gibs_42_reset = reset;
  assign gibs_42_io_cfg_en = cfgRegs_9[44]; // @[CGRA.scala 509:38]
  assign gibs_42_io_cfg_addr = cfgRegs_9[43:32]; // @[CGRA.scala 510:38]
  assign gibs_42_io_cfg_data = cfgRegs_9[31:0]; // @[CGRA.scala 511:38]
  assign gibs_42_io_opinNW_0 = pes_29_io_out_0; // @[CGRA.scala 401:47]
  assign gibs_42_io_opinNE_0 = pes_30_io_out_0; // @[CGRA.scala 400:45]
  assign gibs_42_io_opinSE_0 = pes_38_io_out_0; // @[CGRA.scala 398:41]
  assign gibs_42_io_opinSW_0 = pes_37_io_out_0; // @[CGRA.scala 399:43]
  assign gibs_42_io_itrackW_0 = gibs_41_io_otrackE_0; // @[CGRA.scala 466:16]
  assign gibs_42_io_itrackN_0 = gibs_33_io_otrackS_0; // @[CGRA.scala 436:16]
  assign gibs_42_io_itrackE_0 = gibs_43_io_otrackW_0; // @[CGRA.scala 472:16]
  assign gibs_42_io_itrackS_0 = gibs_51_io_otrackN_0; // @[CGRA.scala 442:16]
  assign gibs_43_clock = clock;
  assign gibs_43_reset = reset;
  assign gibs_43_io_cfg_en = cfgRegs_9[44]; // @[CGRA.scala 509:38]
  assign gibs_43_io_cfg_addr = cfgRegs_9[43:32]; // @[CGRA.scala 510:38]
  assign gibs_43_io_cfg_data = cfgRegs_9[31:0]; // @[CGRA.scala 511:38]
  assign gibs_43_io_opinNW_0 = pes_30_io_out_0; // @[CGRA.scala 401:47]
  assign gibs_43_io_opinNE_0 = pes_31_io_out_0; // @[CGRA.scala 400:45]
  assign gibs_43_io_opinSE_0 = pes_39_io_out_0; // @[CGRA.scala 398:41]
  assign gibs_43_io_opinSW_0 = pes_38_io_out_0; // @[CGRA.scala 399:43]
  assign gibs_43_io_itrackW_0 = gibs_42_io_otrackE_0; // @[CGRA.scala 466:16]
  assign gibs_43_io_itrackN_0 = gibs_34_io_otrackS_0; // @[CGRA.scala 436:16]
  assign gibs_43_io_itrackE_0 = gibs_44_io_otrackW_0; // @[CGRA.scala 472:16]
  assign gibs_43_io_itrackS_0 = gibs_52_io_otrackN_0; // @[CGRA.scala 442:16]
  assign gibs_44_clock = clock;
  assign gibs_44_reset = reset;
  assign gibs_44_io_cfg_en = cfgRegs_9[44]; // @[CGRA.scala 509:38]
  assign gibs_44_io_cfg_addr = cfgRegs_9[43:32]; // @[CGRA.scala 510:38]
  assign gibs_44_io_cfg_data = cfgRegs_9[31:0]; // @[CGRA.scala 511:38]
  assign gibs_44_io_opinNW_0 = pes_31_io_out_0; // @[CGRA.scala 401:47]
  assign gibs_44_io_opinSW_0 = pes_39_io_out_0; // @[CGRA.scala 399:43]
  assign gibs_44_io_itrackW_0 = gibs_43_io_otrackE_0; // @[CGRA.scala 459:16]
  assign gibs_44_io_itrackN_0 = gibs_35_io_otrackS_0; // @[CGRA.scala 436:16]
  assign gibs_44_io_itrackS_0 = gibs_53_io_otrackN_0; // @[CGRA.scala 442:16]
  assign gibs_45_clock = clock;
  assign gibs_45_reset = reset;
  assign gibs_45_io_cfg_en = cfgRegs_11[44]; // @[CGRA.scala 509:38]
  assign gibs_45_io_cfg_addr = cfgRegs_11[43:32]; // @[CGRA.scala 510:38]
  assign gibs_45_io_cfg_data = cfgRegs_11[31:0]; // @[CGRA.scala 511:38]
  assign gibs_45_io_opinNE_0 = pes_32_io_out_0; // @[CGRA.scala 400:45]
  assign gibs_45_io_opinSE_0 = pes_40_io_out_0; // @[CGRA.scala 398:41]
  assign gibs_45_io_itrackN_0 = gibs_36_io_otrackS_0; // @[CGRA.scala 436:16]
  assign gibs_45_io_itrackE_0 = gibs_46_io_otrackW_0; // @[CGRA.scala 451:16]
  assign gibs_45_io_itrackS_0 = gibs_54_io_otrackN_0; // @[CGRA.scala 442:16]
  assign gibs_46_clock = clock;
  assign gibs_46_reset = reset;
  assign gibs_46_io_cfg_en = cfgRegs_11[44]; // @[CGRA.scala 509:38]
  assign gibs_46_io_cfg_addr = cfgRegs_11[43:32]; // @[CGRA.scala 510:38]
  assign gibs_46_io_cfg_data = cfgRegs_11[31:0]; // @[CGRA.scala 511:38]
  assign gibs_46_io_opinNW_0 = pes_32_io_out_0; // @[CGRA.scala 401:47]
  assign gibs_46_io_opinNE_0 = pes_33_io_out_0; // @[CGRA.scala 400:45]
  assign gibs_46_io_opinSE_0 = pes_41_io_out_0; // @[CGRA.scala 398:41]
  assign gibs_46_io_opinSW_0 = pes_40_io_out_0; // @[CGRA.scala 399:43]
  assign gibs_46_io_itrackW_0 = gibs_45_io_otrackE_0; // @[CGRA.scala 466:16]
  assign gibs_46_io_itrackN_0 = gibs_37_io_otrackS_0; // @[CGRA.scala 436:16]
  assign gibs_46_io_itrackE_0 = gibs_47_io_otrackW_0; // @[CGRA.scala 472:16]
  assign gibs_46_io_itrackS_0 = gibs_55_io_otrackN_0; // @[CGRA.scala 442:16]
  assign gibs_47_clock = clock;
  assign gibs_47_reset = reset;
  assign gibs_47_io_cfg_en = cfgRegs_11[44]; // @[CGRA.scala 509:38]
  assign gibs_47_io_cfg_addr = cfgRegs_11[43:32]; // @[CGRA.scala 510:38]
  assign gibs_47_io_cfg_data = cfgRegs_11[31:0]; // @[CGRA.scala 511:38]
  assign gibs_47_io_opinNW_0 = pes_33_io_out_0; // @[CGRA.scala 401:47]
  assign gibs_47_io_opinNE_0 = pes_34_io_out_0; // @[CGRA.scala 400:45]
  assign gibs_47_io_opinSE_0 = pes_42_io_out_0; // @[CGRA.scala 398:41]
  assign gibs_47_io_opinSW_0 = pes_41_io_out_0; // @[CGRA.scala 399:43]
  assign gibs_47_io_itrackW_0 = gibs_46_io_otrackE_0; // @[CGRA.scala 466:16]
  assign gibs_47_io_itrackN_0 = gibs_38_io_otrackS_0; // @[CGRA.scala 436:16]
  assign gibs_47_io_itrackE_0 = gibs_48_io_otrackW_0; // @[CGRA.scala 472:16]
  assign gibs_47_io_itrackS_0 = gibs_56_io_otrackN_0; // @[CGRA.scala 442:16]
  assign gibs_48_clock = clock;
  assign gibs_48_reset = reset;
  assign gibs_48_io_cfg_en = cfgRegs_11[44]; // @[CGRA.scala 509:38]
  assign gibs_48_io_cfg_addr = cfgRegs_11[43:32]; // @[CGRA.scala 510:38]
  assign gibs_48_io_cfg_data = cfgRegs_11[31:0]; // @[CGRA.scala 511:38]
  assign gibs_48_io_opinNW_0 = pes_34_io_out_0; // @[CGRA.scala 401:47]
  assign gibs_48_io_opinNE_0 = pes_35_io_out_0; // @[CGRA.scala 400:45]
  assign gibs_48_io_opinSE_0 = pes_43_io_out_0; // @[CGRA.scala 398:41]
  assign gibs_48_io_opinSW_0 = pes_42_io_out_0; // @[CGRA.scala 399:43]
  assign gibs_48_io_itrackW_0 = gibs_47_io_otrackE_0; // @[CGRA.scala 466:16]
  assign gibs_48_io_itrackN_0 = gibs_39_io_otrackS_0; // @[CGRA.scala 436:16]
  assign gibs_48_io_itrackE_0 = gibs_49_io_otrackW_0; // @[CGRA.scala 472:16]
  assign gibs_48_io_itrackS_0 = gibs_57_io_otrackN_0; // @[CGRA.scala 442:16]
  assign gibs_49_clock = clock;
  assign gibs_49_reset = reset;
  assign gibs_49_io_cfg_en = cfgRegs_11[44]; // @[CGRA.scala 509:38]
  assign gibs_49_io_cfg_addr = cfgRegs_11[43:32]; // @[CGRA.scala 510:38]
  assign gibs_49_io_cfg_data = cfgRegs_11[31:0]; // @[CGRA.scala 511:38]
  assign gibs_49_io_opinNW_0 = pes_35_io_out_0; // @[CGRA.scala 401:47]
  assign gibs_49_io_opinNE_0 = pes_36_io_out_0; // @[CGRA.scala 400:45]
  assign gibs_49_io_opinSE_0 = pes_44_io_out_0; // @[CGRA.scala 398:41]
  assign gibs_49_io_opinSW_0 = pes_43_io_out_0; // @[CGRA.scala 399:43]
  assign gibs_49_io_itrackW_0 = gibs_48_io_otrackE_0; // @[CGRA.scala 466:16]
  assign gibs_49_io_itrackN_0 = gibs_40_io_otrackS_0; // @[CGRA.scala 436:16]
  assign gibs_49_io_itrackE_0 = gibs_50_io_otrackW_0; // @[CGRA.scala 472:16]
  assign gibs_49_io_itrackS_0 = gibs_58_io_otrackN_0; // @[CGRA.scala 442:16]
  assign gibs_50_clock = clock;
  assign gibs_50_reset = reset;
  assign gibs_50_io_cfg_en = cfgRegs_11[44]; // @[CGRA.scala 509:38]
  assign gibs_50_io_cfg_addr = cfgRegs_11[43:32]; // @[CGRA.scala 510:38]
  assign gibs_50_io_cfg_data = cfgRegs_11[31:0]; // @[CGRA.scala 511:38]
  assign gibs_50_io_opinNW_0 = pes_36_io_out_0; // @[CGRA.scala 401:47]
  assign gibs_50_io_opinNE_0 = pes_37_io_out_0; // @[CGRA.scala 400:45]
  assign gibs_50_io_opinSE_0 = pes_45_io_out_0; // @[CGRA.scala 398:41]
  assign gibs_50_io_opinSW_0 = pes_44_io_out_0; // @[CGRA.scala 399:43]
  assign gibs_50_io_itrackW_0 = gibs_49_io_otrackE_0; // @[CGRA.scala 466:16]
  assign gibs_50_io_itrackN_0 = gibs_41_io_otrackS_0; // @[CGRA.scala 436:16]
  assign gibs_50_io_itrackE_0 = gibs_51_io_otrackW_0; // @[CGRA.scala 472:16]
  assign gibs_50_io_itrackS_0 = gibs_59_io_otrackN_0; // @[CGRA.scala 442:16]
  assign gibs_51_clock = clock;
  assign gibs_51_reset = reset;
  assign gibs_51_io_cfg_en = cfgRegs_11[44]; // @[CGRA.scala 509:38]
  assign gibs_51_io_cfg_addr = cfgRegs_11[43:32]; // @[CGRA.scala 510:38]
  assign gibs_51_io_cfg_data = cfgRegs_11[31:0]; // @[CGRA.scala 511:38]
  assign gibs_51_io_opinNW_0 = pes_37_io_out_0; // @[CGRA.scala 401:47]
  assign gibs_51_io_opinNE_0 = pes_38_io_out_0; // @[CGRA.scala 400:45]
  assign gibs_51_io_opinSE_0 = pes_46_io_out_0; // @[CGRA.scala 398:41]
  assign gibs_51_io_opinSW_0 = pes_45_io_out_0; // @[CGRA.scala 399:43]
  assign gibs_51_io_itrackW_0 = gibs_50_io_otrackE_0; // @[CGRA.scala 466:16]
  assign gibs_51_io_itrackN_0 = gibs_42_io_otrackS_0; // @[CGRA.scala 436:16]
  assign gibs_51_io_itrackE_0 = gibs_52_io_otrackW_0; // @[CGRA.scala 472:16]
  assign gibs_51_io_itrackS_0 = gibs_60_io_otrackN_0; // @[CGRA.scala 442:16]
  assign gibs_52_clock = clock;
  assign gibs_52_reset = reset;
  assign gibs_52_io_cfg_en = cfgRegs_11[44]; // @[CGRA.scala 509:38]
  assign gibs_52_io_cfg_addr = cfgRegs_11[43:32]; // @[CGRA.scala 510:38]
  assign gibs_52_io_cfg_data = cfgRegs_11[31:0]; // @[CGRA.scala 511:38]
  assign gibs_52_io_opinNW_0 = pes_38_io_out_0; // @[CGRA.scala 401:47]
  assign gibs_52_io_opinNE_0 = pes_39_io_out_0; // @[CGRA.scala 400:45]
  assign gibs_52_io_opinSE_0 = pes_47_io_out_0; // @[CGRA.scala 398:41]
  assign gibs_52_io_opinSW_0 = pes_46_io_out_0; // @[CGRA.scala 399:43]
  assign gibs_52_io_itrackW_0 = gibs_51_io_otrackE_0; // @[CGRA.scala 466:16]
  assign gibs_52_io_itrackN_0 = gibs_43_io_otrackS_0; // @[CGRA.scala 436:16]
  assign gibs_52_io_itrackE_0 = gibs_53_io_otrackW_0; // @[CGRA.scala 472:16]
  assign gibs_52_io_itrackS_0 = gibs_61_io_otrackN_0; // @[CGRA.scala 442:16]
  assign gibs_53_clock = clock;
  assign gibs_53_reset = reset;
  assign gibs_53_io_cfg_en = cfgRegs_11[44]; // @[CGRA.scala 509:38]
  assign gibs_53_io_cfg_addr = cfgRegs_11[43:32]; // @[CGRA.scala 510:38]
  assign gibs_53_io_cfg_data = cfgRegs_11[31:0]; // @[CGRA.scala 511:38]
  assign gibs_53_io_opinNW_0 = pes_39_io_out_0; // @[CGRA.scala 401:47]
  assign gibs_53_io_opinSW_0 = pes_47_io_out_0; // @[CGRA.scala 399:43]
  assign gibs_53_io_itrackW_0 = gibs_52_io_otrackE_0; // @[CGRA.scala 459:16]
  assign gibs_53_io_itrackN_0 = gibs_44_io_otrackS_0; // @[CGRA.scala 436:16]
  assign gibs_53_io_itrackS_0 = gibs_62_io_otrackN_0; // @[CGRA.scala 442:16]
  assign gibs_54_clock = clock;
  assign gibs_54_reset = reset;
  assign gibs_54_io_cfg_en = cfgRegs_13[44]; // @[CGRA.scala 509:38]
  assign gibs_54_io_cfg_addr = cfgRegs_13[43:32]; // @[CGRA.scala 510:38]
  assign gibs_54_io_cfg_data = cfgRegs_13[31:0]; // @[CGRA.scala 511:38]
  assign gibs_54_io_opinNE_0 = pes_40_io_out_0; // @[CGRA.scala 400:45]
  assign gibs_54_io_opinSE_0 = pes_48_io_out_0; // @[CGRA.scala 398:41]
  assign gibs_54_io_itrackN_0 = gibs_45_io_otrackS_0; // @[CGRA.scala 436:16]
  assign gibs_54_io_itrackE_0 = gibs_55_io_otrackW_0; // @[CGRA.scala 451:16]
  assign gibs_54_io_itrackS_0 = gibs_63_io_otrackN_0; // @[CGRA.scala 442:16]
  assign gibs_55_clock = clock;
  assign gibs_55_reset = reset;
  assign gibs_55_io_cfg_en = cfgRegs_13[44]; // @[CGRA.scala 509:38]
  assign gibs_55_io_cfg_addr = cfgRegs_13[43:32]; // @[CGRA.scala 510:38]
  assign gibs_55_io_cfg_data = cfgRegs_13[31:0]; // @[CGRA.scala 511:38]
  assign gibs_55_io_opinNW_0 = pes_40_io_out_0; // @[CGRA.scala 401:47]
  assign gibs_55_io_opinNE_0 = pes_41_io_out_0; // @[CGRA.scala 400:45]
  assign gibs_55_io_opinSE_0 = pes_49_io_out_0; // @[CGRA.scala 398:41]
  assign gibs_55_io_opinSW_0 = pes_48_io_out_0; // @[CGRA.scala 399:43]
  assign gibs_55_io_itrackW_0 = gibs_54_io_otrackE_0; // @[CGRA.scala 466:16]
  assign gibs_55_io_itrackN_0 = gibs_46_io_otrackS_0; // @[CGRA.scala 436:16]
  assign gibs_55_io_itrackE_0 = gibs_56_io_otrackW_0; // @[CGRA.scala 472:16]
  assign gibs_55_io_itrackS_0 = gibs_64_io_otrackN_0; // @[CGRA.scala 442:16]
  assign gibs_56_clock = clock;
  assign gibs_56_reset = reset;
  assign gibs_56_io_cfg_en = cfgRegs_13[44]; // @[CGRA.scala 509:38]
  assign gibs_56_io_cfg_addr = cfgRegs_13[43:32]; // @[CGRA.scala 510:38]
  assign gibs_56_io_cfg_data = cfgRegs_13[31:0]; // @[CGRA.scala 511:38]
  assign gibs_56_io_opinNW_0 = pes_41_io_out_0; // @[CGRA.scala 401:47]
  assign gibs_56_io_opinNE_0 = pes_42_io_out_0; // @[CGRA.scala 400:45]
  assign gibs_56_io_opinSE_0 = pes_50_io_out_0; // @[CGRA.scala 398:41]
  assign gibs_56_io_opinSW_0 = pes_49_io_out_0; // @[CGRA.scala 399:43]
  assign gibs_56_io_itrackW_0 = gibs_55_io_otrackE_0; // @[CGRA.scala 466:16]
  assign gibs_56_io_itrackN_0 = gibs_47_io_otrackS_0; // @[CGRA.scala 436:16]
  assign gibs_56_io_itrackE_0 = gibs_57_io_otrackW_0; // @[CGRA.scala 472:16]
  assign gibs_56_io_itrackS_0 = gibs_65_io_otrackN_0; // @[CGRA.scala 442:16]
  assign gibs_57_clock = clock;
  assign gibs_57_reset = reset;
  assign gibs_57_io_cfg_en = cfgRegs_13[44]; // @[CGRA.scala 509:38]
  assign gibs_57_io_cfg_addr = cfgRegs_13[43:32]; // @[CGRA.scala 510:38]
  assign gibs_57_io_cfg_data = cfgRegs_13[31:0]; // @[CGRA.scala 511:38]
  assign gibs_57_io_opinNW_0 = pes_42_io_out_0; // @[CGRA.scala 401:47]
  assign gibs_57_io_opinNE_0 = pes_43_io_out_0; // @[CGRA.scala 400:45]
  assign gibs_57_io_opinSE_0 = pes_51_io_out_0; // @[CGRA.scala 398:41]
  assign gibs_57_io_opinSW_0 = pes_50_io_out_0; // @[CGRA.scala 399:43]
  assign gibs_57_io_itrackW_0 = gibs_56_io_otrackE_0; // @[CGRA.scala 466:16]
  assign gibs_57_io_itrackN_0 = gibs_48_io_otrackS_0; // @[CGRA.scala 436:16]
  assign gibs_57_io_itrackE_0 = gibs_58_io_otrackW_0; // @[CGRA.scala 472:16]
  assign gibs_57_io_itrackS_0 = gibs_66_io_otrackN_0; // @[CGRA.scala 442:16]
  assign gibs_58_clock = clock;
  assign gibs_58_reset = reset;
  assign gibs_58_io_cfg_en = cfgRegs_13[44]; // @[CGRA.scala 509:38]
  assign gibs_58_io_cfg_addr = cfgRegs_13[43:32]; // @[CGRA.scala 510:38]
  assign gibs_58_io_cfg_data = cfgRegs_13[31:0]; // @[CGRA.scala 511:38]
  assign gibs_58_io_opinNW_0 = pes_43_io_out_0; // @[CGRA.scala 401:47]
  assign gibs_58_io_opinNE_0 = pes_44_io_out_0; // @[CGRA.scala 400:45]
  assign gibs_58_io_opinSE_0 = pes_52_io_out_0; // @[CGRA.scala 398:41]
  assign gibs_58_io_opinSW_0 = pes_51_io_out_0; // @[CGRA.scala 399:43]
  assign gibs_58_io_itrackW_0 = gibs_57_io_otrackE_0; // @[CGRA.scala 466:16]
  assign gibs_58_io_itrackN_0 = gibs_49_io_otrackS_0; // @[CGRA.scala 436:16]
  assign gibs_58_io_itrackE_0 = gibs_59_io_otrackW_0; // @[CGRA.scala 472:16]
  assign gibs_58_io_itrackS_0 = gibs_67_io_otrackN_0; // @[CGRA.scala 442:16]
  assign gibs_59_clock = clock;
  assign gibs_59_reset = reset;
  assign gibs_59_io_cfg_en = cfgRegs_13[44]; // @[CGRA.scala 509:38]
  assign gibs_59_io_cfg_addr = cfgRegs_13[43:32]; // @[CGRA.scala 510:38]
  assign gibs_59_io_cfg_data = cfgRegs_13[31:0]; // @[CGRA.scala 511:38]
  assign gibs_59_io_opinNW_0 = pes_44_io_out_0; // @[CGRA.scala 401:47]
  assign gibs_59_io_opinNE_0 = pes_45_io_out_0; // @[CGRA.scala 400:45]
  assign gibs_59_io_opinSE_0 = pes_53_io_out_0; // @[CGRA.scala 398:41]
  assign gibs_59_io_opinSW_0 = pes_52_io_out_0; // @[CGRA.scala 399:43]
  assign gibs_59_io_itrackW_0 = gibs_58_io_otrackE_0; // @[CGRA.scala 466:16]
  assign gibs_59_io_itrackN_0 = gibs_50_io_otrackS_0; // @[CGRA.scala 436:16]
  assign gibs_59_io_itrackE_0 = gibs_60_io_otrackW_0; // @[CGRA.scala 472:16]
  assign gibs_59_io_itrackS_0 = gibs_68_io_otrackN_0; // @[CGRA.scala 442:16]
  assign gibs_60_clock = clock;
  assign gibs_60_reset = reset;
  assign gibs_60_io_cfg_en = cfgRegs_13[44]; // @[CGRA.scala 509:38]
  assign gibs_60_io_cfg_addr = cfgRegs_13[43:32]; // @[CGRA.scala 510:38]
  assign gibs_60_io_cfg_data = cfgRegs_13[31:0]; // @[CGRA.scala 511:38]
  assign gibs_60_io_opinNW_0 = pes_45_io_out_0; // @[CGRA.scala 401:47]
  assign gibs_60_io_opinNE_0 = pes_46_io_out_0; // @[CGRA.scala 400:45]
  assign gibs_60_io_opinSE_0 = pes_54_io_out_0; // @[CGRA.scala 398:41]
  assign gibs_60_io_opinSW_0 = pes_53_io_out_0; // @[CGRA.scala 399:43]
  assign gibs_60_io_itrackW_0 = gibs_59_io_otrackE_0; // @[CGRA.scala 466:16]
  assign gibs_60_io_itrackN_0 = gibs_51_io_otrackS_0; // @[CGRA.scala 436:16]
  assign gibs_60_io_itrackE_0 = gibs_61_io_otrackW_0; // @[CGRA.scala 472:16]
  assign gibs_60_io_itrackS_0 = gibs_69_io_otrackN_0; // @[CGRA.scala 442:16]
  assign gibs_61_clock = clock;
  assign gibs_61_reset = reset;
  assign gibs_61_io_cfg_en = cfgRegs_13[44]; // @[CGRA.scala 509:38]
  assign gibs_61_io_cfg_addr = cfgRegs_13[43:32]; // @[CGRA.scala 510:38]
  assign gibs_61_io_cfg_data = cfgRegs_13[31:0]; // @[CGRA.scala 511:38]
  assign gibs_61_io_opinNW_0 = pes_46_io_out_0; // @[CGRA.scala 401:47]
  assign gibs_61_io_opinNE_0 = pes_47_io_out_0; // @[CGRA.scala 400:45]
  assign gibs_61_io_opinSE_0 = pes_55_io_out_0; // @[CGRA.scala 398:41]
  assign gibs_61_io_opinSW_0 = pes_54_io_out_0; // @[CGRA.scala 399:43]
  assign gibs_61_io_itrackW_0 = gibs_60_io_otrackE_0; // @[CGRA.scala 466:16]
  assign gibs_61_io_itrackN_0 = gibs_52_io_otrackS_0; // @[CGRA.scala 436:16]
  assign gibs_61_io_itrackE_0 = gibs_62_io_otrackW_0; // @[CGRA.scala 472:16]
  assign gibs_61_io_itrackS_0 = gibs_70_io_otrackN_0; // @[CGRA.scala 442:16]
  assign gibs_62_clock = clock;
  assign gibs_62_reset = reset;
  assign gibs_62_io_cfg_en = cfgRegs_13[44]; // @[CGRA.scala 509:38]
  assign gibs_62_io_cfg_addr = cfgRegs_13[43:32]; // @[CGRA.scala 510:38]
  assign gibs_62_io_cfg_data = cfgRegs_13[31:0]; // @[CGRA.scala 511:38]
  assign gibs_62_io_opinNW_0 = pes_47_io_out_0; // @[CGRA.scala 401:47]
  assign gibs_62_io_opinSW_0 = pes_55_io_out_0; // @[CGRA.scala 399:43]
  assign gibs_62_io_itrackW_0 = gibs_61_io_otrackE_0; // @[CGRA.scala 459:16]
  assign gibs_62_io_itrackN_0 = gibs_53_io_otrackS_0; // @[CGRA.scala 436:16]
  assign gibs_62_io_itrackS_0 = gibs_71_io_otrackN_0; // @[CGRA.scala 442:16]
  assign gibs_63_clock = clock;
  assign gibs_63_reset = reset;
  assign gibs_63_io_cfg_en = cfgRegs_15[44]; // @[CGRA.scala 509:38]
  assign gibs_63_io_cfg_addr = cfgRegs_15[43:32]; // @[CGRA.scala 510:38]
  assign gibs_63_io_cfg_data = cfgRegs_15[31:0]; // @[CGRA.scala 511:38]
  assign gibs_63_io_opinNE_0 = pes_48_io_out_0; // @[CGRA.scala 400:45]
  assign gibs_63_io_opinSE_0 = pes_56_io_out_0; // @[CGRA.scala 398:41]
  assign gibs_63_io_itrackN_0 = gibs_54_io_otrackS_0; // @[CGRA.scala 436:16]
  assign gibs_63_io_itrackE_0 = gibs_64_io_otrackW_0; // @[CGRA.scala 451:16]
  assign gibs_63_io_itrackS_0 = gibs_72_io_otrackN_0; // @[CGRA.scala 442:16]
  assign gibs_64_clock = clock;
  assign gibs_64_reset = reset;
  assign gibs_64_io_cfg_en = cfgRegs_15[44]; // @[CGRA.scala 509:38]
  assign gibs_64_io_cfg_addr = cfgRegs_15[43:32]; // @[CGRA.scala 510:38]
  assign gibs_64_io_cfg_data = cfgRegs_15[31:0]; // @[CGRA.scala 511:38]
  assign gibs_64_io_opinNW_0 = pes_48_io_out_0; // @[CGRA.scala 401:47]
  assign gibs_64_io_opinNE_0 = pes_49_io_out_0; // @[CGRA.scala 400:45]
  assign gibs_64_io_opinSE_0 = pes_57_io_out_0; // @[CGRA.scala 398:41]
  assign gibs_64_io_opinSW_0 = pes_56_io_out_0; // @[CGRA.scala 399:43]
  assign gibs_64_io_itrackW_0 = gibs_63_io_otrackE_0; // @[CGRA.scala 466:16]
  assign gibs_64_io_itrackN_0 = gibs_55_io_otrackS_0; // @[CGRA.scala 436:16]
  assign gibs_64_io_itrackE_0 = gibs_65_io_otrackW_0; // @[CGRA.scala 472:16]
  assign gibs_64_io_itrackS_0 = gibs_73_io_otrackN_0; // @[CGRA.scala 442:16]
  assign gibs_65_clock = clock;
  assign gibs_65_reset = reset;
  assign gibs_65_io_cfg_en = cfgRegs_15[44]; // @[CGRA.scala 509:38]
  assign gibs_65_io_cfg_addr = cfgRegs_15[43:32]; // @[CGRA.scala 510:38]
  assign gibs_65_io_cfg_data = cfgRegs_15[31:0]; // @[CGRA.scala 511:38]
  assign gibs_65_io_opinNW_0 = pes_49_io_out_0; // @[CGRA.scala 401:47]
  assign gibs_65_io_opinNE_0 = pes_50_io_out_0; // @[CGRA.scala 400:45]
  assign gibs_65_io_opinSE_0 = pes_58_io_out_0; // @[CGRA.scala 398:41]
  assign gibs_65_io_opinSW_0 = pes_57_io_out_0; // @[CGRA.scala 399:43]
  assign gibs_65_io_itrackW_0 = gibs_64_io_otrackE_0; // @[CGRA.scala 466:16]
  assign gibs_65_io_itrackN_0 = gibs_56_io_otrackS_0; // @[CGRA.scala 436:16]
  assign gibs_65_io_itrackE_0 = gibs_66_io_otrackW_0; // @[CGRA.scala 472:16]
  assign gibs_65_io_itrackS_0 = gibs_74_io_otrackN_0; // @[CGRA.scala 442:16]
  assign gibs_66_clock = clock;
  assign gibs_66_reset = reset;
  assign gibs_66_io_cfg_en = cfgRegs_15[44]; // @[CGRA.scala 509:38]
  assign gibs_66_io_cfg_addr = cfgRegs_15[43:32]; // @[CGRA.scala 510:38]
  assign gibs_66_io_cfg_data = cfgRegs_15[31:0]; // @[CGRA.scala 511:38]
  assign gibs_66_io_opinNW_0 = pes_50_io_out_0; // @[CGRA.scala 401:47]
  assign gibs_66_io_opinNE_0 = pes_51_io_out_0; // @[CGRA.scala 400:45]
  assign gibs_66_io_opinSE_0 = pes_59_io_out_0; // @[CGRA.scala 398:41]
  assign gibs_66_io_opinSW_0 = pes_58_io_out_0; // @[CGRA.scala 399:43]
  assign gibs_66_io_itrackW_0 = gibs_65_io_otrackE_0; // @[CGRA.scala 466:16]
  assign gibs_66_io_itrackN_0 = gibs_57_io_otrackS_0; // @[CGRA.scala 436:16]
  assign gibs_66_io_itrackE_0 = gibs_67_io_otrackW_0; // @[CGRA.scala 472:16]
  assign gibs_66_io_itrackS_0 = gibs_75_io_otrackN_0; // @[CGRA.scala 442:16]
  assign gibs_67_clock = clock;
  assign gibs_67_reset = reset;
  assign gibs_67_io_cfg_en = cfgRegs_15[44]; // @[CGRA.scala 509:38]
  assign gibs_67_io_cfg_addr = cfgRegs_15[43:32]; // @[CGRA.scala 510:38]
  assign gibs_67_io_cfg_data = cfgRegs_15[31:0]; // @[CGRA.scala 511:38]
  assign gibs_67_io_opinNW_0 = pes_51_io_out_0; // @[CGRA.scala 401:47]
  assign gibs_67_io_opinNE_0 = pes_52_io_out_0; // @[CGRA.scala 400:45]
  assign gibs_67_io_opinSE_0 = pes_60_io_out_0; // @[CGRA.scala 398:41]
  assign gibs_67_io_opinSW_0 = pes_59_io_out_0; // @[CGRA.scala 399:43]
  assign gibs_67_io_itrackW_0 = gibs_66_io_otrackE_0; // @[CGRA.scala 466:16]
  assign gibs_67_io_itrackN_0 = gibs_58_io_otrackS_0; // @[CGRA.scala 436:16]
  assign gibs_67_io_itrackE_0 = gibs_68_io_otrackW_0; // @[CGRA.scala 472:16]
  assign gibs_67_io_itrackS_0 = gibs_76_io_otrackN_0; // @[CGRA.scala 442:16]
  assign gibs_68_clock = clock;
  assign gibs_68_reset = reset;
  assign gibs_68_io_cfg_en = cfgRegs_15[44]; // @[CGRA.scala 509:38]
  assign gibs_68_io_cfg_addr = cfgRegs_15[43:32]; // @[CGRA.scala 510:38]
  assign gibs_68_io_cfg_data = cfgRegs_15[31:0]; // @[CGRA.scala 511:38]
  assign gibs_68_io_opinNW_0 = pes_52_io_out_0; // @[CGRA.scala 401:47]
  assign gibs_68_io_opinNE_0 = pes_53_io_out_0; // @[CGRA.scala 400:45]
  assign gibs_68_io_opinSE_0 = pes_61_io_out_0; // @[CGRA.scala 398:41]
  assign gibs_68_io_opinSW_0 = pes_60_io_out_0; // @[CGRA.scala 399:43]
  assign gibs_68_io_itrackW_0 = gibs_67_io_otrackE_0; // @[CGRA.scala 466:16]
  assign gibs_68_io_itrackN_0 = gibs_59_io_otrackS_0; // @[CGRA.scala 436:16]
  assign gibs_68_io_itrackE_0 = gibs_69_io_otrackW_0; // @[CGRA.scala 472:16]
  assign gibs_68_io_itrackS_0 = gibs_77_io_otrackN_0; // @[CGRA.scala 442:16]
  assign gibs_69_clock = clock;
  assign gibs_69_reset = reset;
  assign gibs_69_io_cfg_en = cfgRegs_15[44]; // @[CGRA.scala 509:38]
  assign gibs_69_io_cfg_addr = cfgRegs_15[43:32]; // @[CGRA.scala 510:38]
  assign gibs_69_io_cfg_data = cfgRegs_15[31:0]; // @[CGRA.scala 511:38]
  assign gibs_69_io_opinNW_0 = pes_53_io_out_0; // @[CGRA.scala 401:47]
  assign gibs_69_io_opinNE_0 = pes_54_io_out_0; // @[CGRA.scala 400:45]
  assign gibs_69_io_opinSE_0 = pes_62_io_out_0; // @[CGRA.scala 398:41]
  assign gibs_69_io_opinSW_0 = pes_61_io_out_0; // @[CGRA.scala 399:43]
  assign gibs_69_io_itrackW_0 = gibs_68_io_otrackE_0; // @[CGRA.scala 466:16]
  assign gibs_69_io_itrackN_0 = gibs_60_io_otrackS_0; // @[CGRA.scala 436:16]
  assign gibs_69_io_itrackE_0 = gibs_70_io_otrackW_0; // @[CGRA.scala 472:16]
  assign gibs_69_io_itrackS_0 = gibs_78_io_otrackN_0; // @[CGRA.scala 442:16]
  assign gibs_70_clock = clock;
  assign gibs_70_reset = reset;
  assign gibs_70_io_cfg_en = cfgRegs_15[44]; // @[CGRA.scala 509:38]
  assign gibs_70_io_cfg_addr = cfgRegs_15[43:32]; // @[CGRA.scala 510:38]
  assign gibs_70_io_cfg_data = cfgRegs_15[31:0]; // @[CGRA.scala 511:38]
  assign gibs_70_io_opinNW_0 = pes_54_io_out_0; // @[CGRA.scala 401:47]
  assign gibs_70_io_opinNE_0 = pes_55_io_out_0; // @[CGRA.scala 400:45]
  assign gibs_70_io_opinSE_0 = pes_63_io_out_0; // @[CGRA.scala 398:41]
  assign gibs_70_io_opinSW_0 = pes_62_io_out_0; // @[CGRA.scala 399:43]
  assign gibs_70_io_itrackW_0 = gibs_69_io_otrackE_0; // @[CGRA.scala 466:16]
  assign gibs_70_io_itrackN_0 = gibs_61_io_otrackS_0; // @[CGRA.scala 436:16]
  assign gibs_70_io_itrackE_0 = gibs_71_io_otrackW_0; // @[CGRA.scala 472:16]
  assign gibs_70_io_itrackS_0 = gibs_79_io_otrackN_0; // @[CGRA.scala 442:16]
  assign gibs_71_clock = clock;
  assign gibs_71_reset = reset;
  assign gibs_71_io_cfg_en = cfgRegs_15[44]; // @[CGRA.scala 509:38]
  assign gibs_71_io_cfg_addr = cfgRegs_15[43:32]; // @[CGRA.scala 510:38]
  assign gibs_71_io_cfg_data = cfgRegs_15[31:0]; // @[CGRA.scala 511:38]
  assign gibs_71_io_opinNW_0 = pes_55_io_out_0; // @[CGRA.scala 401:47]
  assign gibs_71_io_opinSW_0 = pes_63_io_out_0; // @[CGRA.scala 399:43]
  assign gibs_71_io_itrackW_0 = gibs_70_io_otrackE_0; // @[CGRA.scala 459:16]
  assign gibs_71_io_itrackN_0 = gibs_62_io_otrackS_0; // @[CGRA.scala 436:16]
  assign gibs_71_io_itrackS_0 = gibs_80_io_otrackN_0; // @[CGRA.scala 442:16]
  assign gibs_72_clock = clock;
  assign gibs_72_reset = reset;
  assign gibs_72_io_cfg_en = cfgRegs_17[44]; // @[CGRA.scala 509:38]
  assign gibs_72_io_cfg_addr = cfgRegs_17[43:32]; // @[CGRA.scala 510:38]
  assign gibs_72_io_cfg_data = cfgRegs_17[31:0]; // @[CGRA.scala 511:38]
  assign gibs_72_io_opinNE_0 = pes_56_io_out_0; // @[CGRA.scala 400:45]
  assign gibs_72_io_opinSE_0 = ibs_8_io_out_0; // @[CGRA.scala 334:35]
  assign gibs_72_io_itrackN_0 = gibs_63_io_otrackS_0; // @[CGRA.scala 429:16]
  assign gibs_72_io_itrackE_0 = gibs_73_io_otrackW_0; // @[CGRA.scala 451:16]
  assign gibs_73_clock = clock;
  assign gibs_73_reset = reset;
  assign gibs_73_io_cfg_en = cfgRegs_17[44]; // @[CGRA.scala 509:38]
  assign gibs_73_io_cfg_addr = cfgRegs_17[43:32]; // @[CGRA.scala 510:38]
  assign gibs_73_io_cfg_data = cfgRegs_17[31:0]; // @[CGRA.scala 511:38]
  assign gibs_73_io_opinNW_0 = pes_56_io_out_0; // @[CGRA.scala 401:47]
  assign gibs_73_io_opinNE_0 = pes_57_io_out_0; // @[CGRA.scala 400:45]
  assign gibs_73_io_opinSE_0 = ibs_9_io_out_0; // @[CGRA.scala 334:35]
  assign gibs_73_io_opinSW_0 = ibs_8_io_out_0; // @[CGRA.scala 335:37]
  assign gibs_73_io_itrackW_0 = gibs_72_io_otrackE_0; // @[CGRA.scala 466:16]
  assign gibs_73_io_itrackN_0 = gibs_64_io_otrackS_0; // @[CGRA.scala 429:16]
  assign gibs_73_io_itrackE_0 = gibs_74_io_otrackW_0; // @[CGRA.scala 472:16]
  assign gibs_74_clock = clock;
  assign gibs_74_reset = reset;
  assign gibs_74_io_cfg_en = cfgRegs_17[44]; // @[CGRA.scala 509:38]
  assign gibs_74_io_cfg_addr = cfgRegs_17[43:32]; // @[CGRA.scala 510:38]
  assign gibs_74_io_cfg_data = cfgRegs_17[31:0]; // @[CGRA.scala 511:38]
  assign gibs_74_io_opinNW_0 = pes_57_io_out_0; // @[CGRA.scala 401:47]
  assign gibs_74_io_opinNE_0 = pes_58_io_out_0; // @[CGRA.scala 400:45]
  assign gibs_74_io_opinSE_0 = ibs_10_io_out_0; // @[CGRA.scala 334:35]
  assign gibs_74_io_opinSW_0 = ibs_9_io_out_0; // @[CGRA.scala 335:37]
  assign gibs_74_io_itrackW_0 = gibs_73_io_otrackE_0; // @[CGRA.scala 466:16]
  assign gibs_74_io_itrackN_0 = gibs_65_io_otrackS_0; // @[CGRA.scala 429:16]
  assign gibs_74_io_itrackE_0 = gibs_75_io_otrackW_0; // @[CGRA.scala 472:16]
  assign gibs_75_clock = clock;
  assign gibs_75_reset = reset;
  assign gibs_75_io_cfg_en = cfgRegs_17[44]; // @[CGRA.scala 509:38]
  assign gibs_75_io_cfg_addr = cfgRegs_17[43:32]; // @[CGRA.scala 510:38]
  assign gibs_75_io_cfg_data = cfgRegs_17[31:0]; // @[CGRA.scala 511:38]
  assign gibs_75_io_opinNW_0 = pes_58_io_out_0; // @[CGRA.scala 401:47]
  assign gibs_75_io_opinNE_0 = pes_59_io_out_0; // @[CGRA.scala 400:45]
  assign gibs_75_io_opinSE_0 = ibs_11_io_out_0; // @[CGRA.scala 334:35]
  assign gibs_75_io_opinSW_0 = ibs_10_io_out_0; // @[CGRA.scala 335:37]
  assign gibs_75_io_itrackW_0 = gibs_74_io_otrackE_0; // @[CGRA.scala 466:16]
  assign gibs_75_io_itrackN_0 = gibs_66_io_otrackS_0; // @[CGRA.scala 429:16]
  assign gibs_75_io_itrackE_0 = gibs_76_io_otrackW_0; // @[CGRA.scala 472:16]
  assign gibs_76_clock = clock;
  assign gibs_76_reset = reset;
  assign gibs_76_io_cfg_en = cfgRegs_17[44]; // @[CGRA.scala 509:38]
  assign gibs_76_io_cfg_addr = cfgRegs_17[43:32]; // @[CGRA.scala 510:38]
  assign gibs_76_io_cfg_data = cfgRegs_17[31:0]; // @[CGRA.scala 511:38]
  assign gibs_76_io_opinNW_0 = pes_59_io_out_0; // @[CGRA.scala 401:47]
  assign gibs_76_io_opinNE_0 = pes_60_io_out_0; // @[CGRA.scala 400:45]
  assign gibs_76_io_opinSE_0 = ibs_12_io_out_0; // @[CGRA.scala 334:35]
  assign gibs_76_io_opinSW_0 = ibs_11_io_out_0; // @[CGRA.scala 335:37]
  assign gibs_76_io_itrackW_0 = gibs_75_io_otrackE_0; // @[CGRA.scala 466:16]
  assign gibs_76_io_itrackN_0 = gibs_67_io_otrackS_0; // @[CGRA.scala 429:16]
  assign gibs_76_io_itrackE_0 = gibs_77_io_otrackW_0; // @[CGRA.scala 472:16]
  assign gibs_77_clock = clock;
  assign gibs_77_reset = reset;
  assign gibs_77_io_cfg_en = cfgRegs_17[44]; // @[CGRA.scala 509:38]
  assign gibs_77_io_cfg_addr = cfgRegs_17[43:32]; // @[CGRA.scala 510:38]
  assign gibs_77_io_cfg_data = cfgRegs_17[31:0]; // @[CGRA.scala 511:38]
  assign gibs_77_io_opinNW_0 = pes_60_io_out_0; // @[CGRA.scala 401:47]
  assign gibs_77_io_opinNE_0 = pes_61_io_out_0; // @[CGRA.scala 400:45]
  assign gibs_77_io_opinSE_0 = ibs_13_io_out_0; // @[CGRA.scala 334:35]
  assign gibs_77_io_opinSW_0 = ibs_12_io_out_0; // @[CGRA.scala 335:37]
  assign gibs_77_io_itrackW_0 = gibs_76_io_otrackE_0; // @[CGRA.scala 466:16]
  assign gibs_77_io_itrackN_0 = gibs_68_io_otrackS_0; // @[CGRA.scala 429:16]
  assign gibs_77_io_itrackE_0 = gibs_78_io_otrackW_0; // @[CGRA.scala 472:16]
  assign gibs_78_clock = clock;
  assign gibs_78_reset = reset;
  assign gibs_78_io_cfg_en = cfgRegs_17[44]; // @[CGRA.scala 509:38]
  assign gibs_78_io_cfg_addr = cfgRegs_17[43:32]; // @[CGRA.scala 510:38]
  assign gibs_78_io_cfg_data = cfgRegs_17[31:0]; // @[CGRA.scala 511:38]
  assign gibs_78_io_opinNW_0 = pes_61_io_out_0; // @[CGRA.scala 401:47]
  assign gibs_78_io_opinNE_0 = pes_62_io_out_0; // @[CGRA.scala 400:45]
  assign gibs_78_io_opinSE_0 = ibs_14_io_out_0; // @[CGRA.scala 334:35]
  assign gibs_78_io_opinSW_0 = ibs_13_io_out_0; // @[CGRA.scala 335:37]
  assign gibs_78_io_itrackW_0 = gibs_77_io_otrackE_0; // @[CGRA.scala 466:16]
  assign gibs_78_io_itrackN_0 = gibs_69_io_otrackS_0; // @[CGRA.scala 429:16]
  assign gibs_78_io_itrackE_0 = gibs_79_io_otrackW_0; // @[CGRA.scala 472:16]
  assign gibs_79_clock = clock;
  assign gibs_79_reset = reset;
  assign gibs_79_io_cfg_en = cfgRegs_17[44]; // @[CGRA.scala 509:38]
  assign gibs_79_io_cfg_addr = cfgRegs_17[43:32]; // @[CGRA.scala 510:38]
  assign gibs_79_io_cfg_data = cfgRegs_17[31:0]; // @[CGRA.scala 511:38]
  assign gibs_79_io_opinNW_0 = pes_62_io_out_0; // @[CGRA.scala 401:47]
  assign gibs_79_io_opinNE_0 = pes_63_io_out_0; // @[CGRA.scala 400:45]
  assign gibs_79_io_opinSE_0 = ibs_15_io_out_0; // @[CGRA.scala 334:35]
  assign gibs_79_io_opinSW_0 = ibs_14_io_out_0; // @[CGRA.scala 335:37]
  assign gibs_79_io_itrackW_0 = gibs_78_io_otrackE_0; // @[CGRA.scala 466:16]
  assign gibs_79_io_itrackN_0 = gibs_70_io_otrackS_0; // @[CGRA.scala 429:16]
  assign gibs_79_io_itrackE_0 = gibs_80_io_otrackW_0; // @[CGRA.scala 472:16]
  assign gibs_80_clock = clock;
  assign gibs_80_reset = reset;
  assign gibs_80_io_cfg_en = cfgRegs_17[44]; // @[CGRA.scala 509:38]
  assign gibs_80_io_cfg_addr = cfgRegs_17[43:32]; // @[CGRA.scala 510:38]
  assign gibs_80_io_cfg_data = cfgRegs_17[31:0]; // @[CGRA.scala 511:38]
  assign gibs_80_io_opinNW_0 = pes_63_io_out_0; // @[CGRA.scala 401:47]
  assign gibs_80_io_opinSW_0 = ibs_15_io_out_0; // @[CGRA.scala 335:37]
  assign gibs_80_io_itrackW_0 = gibs_79_io_otrackE_0; // @[CGRA.scala 459:16]
  assign gibs_80_io_itrackN_0 = gibs_71_io_otrackS_0; // @[CGRA.scala 429:16]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  cfgRegs_0 = _RAND_0[44:0];
  _RAND_1 = {2{`RANDOM}};
  cfgRegs_1 = _RAND_1[44:0];
  _RAND_2 = {2{`RANDOM}};
  cfgRegs_2 = _RAND_2[44:0];
  _RAND_3 = {2{`RANDOM}};
  cfgRegs_3 = _RAND_3[44:0];
  _RAND_4 = {2{`RANDOM}};
  cfgRegs_4 = _RAND_4[44:0];
  _RAND_5 = {2{`RANDOM}};
  cfgRegs_5 = _RAND_5[44:0];
  _RAND_6 = {2{`RANDOM}};
  cfgRegs_6 = _RAND_6[44:0];
  _RAND_7 = {2{`RANDOM}};
  cfgRegs_7 = _RAND_7[44:0];
  _RAND_8 = {2{`RANDOM}};
  cfgRegs_8 = _RAND_8[44:0];
  _RAND_9 = {2{`RANDOM}};
  cfgRegs_9 = _RAND_9[44:0];
  _RAND_10 = {2{`RANDOM}};
  cfgRegs_10 = _RAND_10[44:0];
  _RAND_11 = {2{`RANDOM}};
  cfgRegs_11 = _RAND_11[44:0];
  _RAND_12 = {2{`RANDOM}};
  cfgRegs_12 = _RAND_12[44:0];
  _RAND_13 = {2{`RANDOM}};
  cfgRegs_13 = _RAND_13[44:0];
  _RAND_14 = {2{`RANDOM}};
  cfgRegs_14 = _RAND_14[44:0];
  _RAND_15 = {2{`RANDOM}};
  cfgRegs_15 = _RAND_15[44:0];
  _RAND_16 = {2{`RANDOM}};
  cfgRegs_16 = _RAND_16[44:0];
  _RAND_17 = {2{`RANDOM}};
  cfgRegs_17 = _RAND_17[44:0];
  _RAND_18 = {2{`RANDOM}};
  cfgRegs_18 = _RAND_18[44:0];
  _RAND_19 = {2{`RANDOM}};
  cfgRegs_19 = _RAND_19[44:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      cfgRegs_0 <= 45'h0;
    end else begin
      cfgRegs_0 <= _T_2;
    end
    if (reset) begin
      cfgRegs_1 <= 45'h0;
    end else begin
      cfgRegs_1 <= cfgRegs_0;
    end
    if (reset) begin
      cfgRegs_2 <= 45'h0;
    end else begin
      cfgRegs_2 <= cfgRegs_1;
    end
    if (reset) begin
      cfgRegs_3 <= 45'h0;
    end else begin
      cfgRegs_3 <= cfgRegs_2;
    end
    if (reset) begin
      cfgRegs_4 <= 45'h0;
    end else begin
      cfgRegs_4 <= cfgRegs_3;
    end
    if (reset) begin
      cfgRegs_5 <= 45'h0;
    end else begin
      cfgRegs_5 <= cfgRegs_4;
    end
    if (reset) begin
      cfgRegs_6 <= 45'h0;
    end else begin
      cfgRegs_6 <= cfgRegs_5;
    end
    if (reset) begin
      cfgRegs_7 <= 45'h0;
    end else begin
      cfgRegs_7 <= cfgRegs_6;
    end
    if (reset) begin
      cfgRegs_8 <= 45'h0;
    end else begin
      cfgRegs_8 <= cfgRegs_7;
    end
    if (reset) begin
      cfgRegs_9 <= 45'h0;
    end else begin
      cfgRegs_9 <= cfgRegs_8;
    end
    if (reset) begin
      cfgRegs_10 <= 45'h0;
    end else begin
      cfgRegs_10 <= cfgRegs_9;
    end
    if (reset) begin
      cfgRegs_11 <= 45'h0;
    end else begin
      cfgRegs_11 <= cfgRegs_10;
    end
    if (reset) begin
      cfgRegs_12 <= 45'h0;
    end else begin
      cfgRegs_12 <= cfgRegs_11;
    end
    if (reset) begin
      cfgRegs_13 <= 45'h0;
    end else begin
      cfgRegs_13 <= cfgRegs_12;
    end
    if (reset) begin
      cfgRegs_14 <= 45'h0;
    end else begin
      cfgRegs_14 <= cfgRegs_13;
    end
    if (reset) begin
      cfgRegs_15 <= 45'h0;
    end else begin
      cfgRegs_15 <= cfgRegs_14;
    end
    if (reset) begin
      cfgRegs_16 <= 45'h0;
    end else begin
      cfgRegs_16 <= cfgRegs_15;
    end
    if (reset) begin
      cfgRegs_17 <= 45'h0;
    end else begin
      cfgRegs_17 <= cfgRegs_16;
    end
    if (reset) begin
      cfgRegs_18 <= 45'h0;
    end else begin
      cfgRegs_18 <= cfgRegs_17;
    end
    if (reset) begin
      cfgRegs_19 <= 45'h0;
    end else begin
      cfgRegs_19 <= cfgRegs_18;
    end
  end
endmodule
